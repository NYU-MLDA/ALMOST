//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n839_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT78), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT78), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n212_), .A2(new_n205_), .A3(new_n204_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT26), .B(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n215_), .B(new_n218_), .C1(new_n219_), .C2(new_n216_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n208_), .A2(new_n209_), .A3(new_n214_), .A4(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G169gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n212_), .B1(new_n223_), .B2(new_n211_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT79), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G71gat), .B(G99gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n227_), .B(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G127gat), .B(G134gat), .Z(new_n232_));
  XOR2_X1   g031(.A(G113gat), .B(G120gat), .Z(new_n233_));
  XOR2_X1   g032(.A(new_n232_), .B(new_n233_), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G15gat), .B(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT30), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n236_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242_));
  OR2_X1    g041(.A1(G155gat), .A2(G162gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(KEYINPUT3), .Z(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT2), .Z(new_n247_));
  OAI211_X1 g046(.A(new_n242_), .B(new_n243_), .C1(new_n245_), .C2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n244_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT80), .B1(new_n242_), .B2(KEYINPUT1), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(KEYINPUT1), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n243_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n242_), .A2(KEYINPUT80), .A3(KEYINPUT1), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n249_), .B(new_n246_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n254_), .A3(new_n235_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n248_), .A2(new_n254_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n234_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(KEYINPUT92), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT92), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n259_), .A3(new_n234_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n241_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT94), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n264_));
  NAND3_X1  g063(.A1(new_n256_), .A2(new_n234_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n262_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT94), .B1(new_n261_), .B2(new_n268_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT95), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n258_), .A2(new_n260_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(new_n266_), .ZN(new_n274_));
  AOI211_X1 g073(.A(KEYINPUT95), .B(new_n267_), .C1(new_n258_), .C2(new_n260_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n270_), .B(new_n271_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G29gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT0), .ZN(new_n278_));
  INV_X1    g077(.A(G57gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G85gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n274_), .A2(new_n275_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n284_), .A2(new_n281_), .A3(new_n271_), .A4(new_n270_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n240_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G78gat), .B(G106gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT88), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G211gat), .B(G218gat), .Z(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT21), .ZN(new_n293_));
  INV_X1    g092(.A(G197gat), .ZN(new_n294_));
  INV_X1    g093(.A(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT84), .B(G197gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(new_n295_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n295_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(G197gat), .B2(G204gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n292_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT86), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n299_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT83), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n256_), .A2(KEYINPUT29), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT87), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n316_), .A3(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n311_), .A2(new_n313_), .ZN(new_n321_));
  OAI211_X1 g120(.A(KEYINPUT87), .B(new_n318_), .C1(new_n321_), .C2(KEYINPUT83), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n291_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT89), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n291_), .A3(new_n322_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT90), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n320_), .A2(KEYINPUT90), .A3(new_n291_), .A4(new_n322_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(KEYINPUT89), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n256_), .A2(KEYINPUT29), .ZN(new_n331_));
  XOR2_X1   g130(.A(G22gat), .B(G50gat), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT82), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n331_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT81), .B(KEYINPUT28), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n222_), .B(KEYINPUT91), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n213_), .B1(new_n219_), .B2(new_n215_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n338_), .A2(new_n224_), .B1(new_n207_), .B2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(new_n310_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n310_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT20), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n311_), .A2(new_n226_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n345_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n340_), .A2(new_n310_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n347_), .A2(KEYINPUT20), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT18), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G64gat), .ZN(new_n354_));
  INV_X1    g153(.A(G92gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n351_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT27), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n351_), .A2(new_n357_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(new_n359_), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n362_));
  NAND3_X1  g161(.A1(new_n347_), .A2(new_n349_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n345_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n341_), .A2(KEYINPUT20), .A3(new_n348_), .A4(new_n342_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n357_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n358_), .A2(new_n359_), .B1(new_n361_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n336_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n325_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n370_), .A2(new_n323_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n337_), .A2(new_n368_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT98), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n330_), .B2(new_n336_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT98), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n368_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n288_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n351_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n379_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n356_), .B1(new_n346_), .B2(new_n350_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n360_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n286_), .B2(KEYINPUT33), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT96), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n265_), .A2(new_n266_), .ZN(new_n389_));
  OR3_X1    g188(.A1(new_n261_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n261_), .B2(new_n389_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n281_), .B1(new_n273_), .B2(new_n267_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n387_), .B1(new_n285_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n383_), .B1(new_n386_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n375_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n323_), .B(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n327_), .A2(new_n328_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n369_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n368_), .B(new_n287_), .C1(new_n400_), .C2(new_n371_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n240_), .B1(new_n396_), .B2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n378_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G99gat), .A2(G106gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(G85gat), .A2(G92gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT9), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(KEYINPUT65), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT10), .B(G99gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G106gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G85gat), .A2(G92gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n409_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(new_n410_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT65), .B1(new_n409_), .B2(KEYINPUT9), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n412_), .B(new_n416_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT7), .ZN(new_n422_));
  INV_X1    g221(.A(G99gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n415_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n424_), .A2(new_n406_), .A3(new_n407_), .A4(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n409_), .A2(new_n417_), .A3(KEYINPUT8), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT66), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT66), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n430_), .A3(new_n427_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT8), .ZN(new_n433_));
  INV_X1    g232(.A(new_n404_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT67), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(KEYINPUT6), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n405_), .A2(KEYINPUT67), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n434_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n425_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n405_), .A2(KEYINPUT67), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n435_), .A2(KEYINPUT6), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n404_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n438_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n433_), .B1(new_n445_), .B2(new_n418_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n421_), .B1(new_n432_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n404_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n418_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT8), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n426_), .A2(new_n430_), .A3(new_n427_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n430_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(KEYINPUT68), .A3(new_n421_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G71gat), .B(G78gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(G57gat), .B(G64gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(KEYINPUT11), .B2(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(KEYINPUT11), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT12), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n449_), .A2(new_n458_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n447_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n463_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n463_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n447_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT69), .B1(new_n471_), .B2(new_n464_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT69), .ZN(new_n473_));
  AOI211_X1 g272(.A(new_n473_), .B(KEYINPUT12), .C1(new_n447_), .C2(new_n470_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G230gat), .A2(G233gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n476_), .B(KEYINPUT64), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n469_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n468_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n463_), .B1(new_n457_), .B2(new_n421_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G120gat), .B(G148gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(new_n295_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT5), .B(G176gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n486_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT76), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496_));
  INV_X1    g295(.A(G1gat), .ZN(new_n497_));
  INV_X1    g296(.A(G8gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G1gat), .B(G8gat), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(KEYINPUT75), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT75), .ZN(new_n509_));
  INV_X1    g308(.A(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n502_), .A2(new_n503_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n507_), .B(KEYINPUT15), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n511_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n508_), .A2(new_n512_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n519_), .A2(new_n517_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(G169gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(new_n294_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n495_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n518_), .A2(new_n520_), .A3(KEYINPUT76), .A4(new_n524_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n494_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n403_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT35), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G232gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT70), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT34), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n467_), .A2(new_n507_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n449_), .A2(new_n458_), .A3(new_n514_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n538_), .A2(new_n535_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n539_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G134gat), .B(G162gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  OR4_X1    g346(.A1(KEYINPUT36), .A2(new_n543_), .A3(new_n544_), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n547_), .B(KEYINPUT36), .Z(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT37), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n511_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n463_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n558_));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT72), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n562_), .A2(new_n563_), .A3(KEYINPUT17), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(KEYINPUT17), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n557_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n564_), .B2(new_n557_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT74), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n554_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n534_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n287_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n497_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT38), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n288_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n377_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n376_), .B1(new_n375_), .B2(new_n368_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n396_), .A2(new_n401_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n236_), .B(new_n239_), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n548_), .A2(new_n551_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n532_), .A2(new_n568_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT99), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n497_), .B1(new_n590_), .B2(new_n573_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n576_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n574_), .A2(new_n593_), .A3(new_n575_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT101), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n592_), .B(new_n599_), .C1(new_n594_), .C2(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(G1324gat));
  INV_X1    g400(.A(new_n368_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n572_), .A2(new_n498_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n498_), .B1(new_n590_), .B2(new_n602_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n604_), .A2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n603_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT40), .B(new_n603_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1325gat));
  OAI21_X1  g412(.A(G15gat), .B1(new_n589_), .B2(new_n582_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT102), .Z(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT41), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT41), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n571_), .A2(G15gat), .A3(new_n582_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n589_), .B2(new_n375_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n375_), .A2(G22gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n571_), .B2(new_n622_), .ZN(G1327gat));
  NOR2_X1   g422(.A1(new_n568_), .A2(new_n585_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT104), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n534_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n573_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n532_), .A2(new_n569_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n584_), .B2(new_n554_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n631_), .B(new_n554_), .C1(new_n378_), .C2(new_n402_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT44), .B(new_n630_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n635_), .A2(G29gat), .A3(new_n573_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n632_), .A2(new_n634_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n629_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n628_), .B1(new_n636_), .B2(new_n640_), .ZN(G1328gat));
  OAI21_X1  g440(.A(KEYINPUT43), .B1(new_n403_), .B2(new_n553_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n629_), .B1(new_n642_), .B2(new_n633_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n635_), .B(new_n602_), .C1(new_n643_), .C2(new_n637_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT105), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n640_), .A2(new_n646_), .A3(new_n602_), .A4(new_n635_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n647_), .A3(G36gat), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n368_), .A2(G36gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT106), .B1(new_n626_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n534_), .A2(new_n652_), .A3(new_n625_), .A4(new_n649_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n651_), .A2(KEYINPUT45), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT45), .B1(new_n651_), .B2(new_n653_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n648_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT108), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n648_), .A2(new_n659_), .A3(new_n656_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1329gat));
  NOR3_X1   g462(.A1(new_n626_), .A2(G43gat), .A3(new_n582_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n640_), .A2(new_n240_), .A3(new_n635_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(G43gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g466(.A(new_n375_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n640_), .A2(new_n668_), .A3(new_n635_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G50gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n375_), .A2(G50gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT109), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n626_), .B2(new_n672_), .ZN(G1331gat));
  NAND4_X1  g472(.A1(new_n586_), .A2(new_n568_), .A3(new_n531_), .A4(new_n494_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(new_n279_), .A3(new_n287_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n584_), .A2(new_n531_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT110), .ZN(new_n677_));
  INV_X1    g476(.A(new_n494_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n570_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n279_), .B1(new_n680_), .B2(new_n287_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT111), .B(new_n279_), .C1(new_n680_), .C2(new_n287_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n675_), .B1(new_n683_), .B2(new_n684_), .ZN(G1332gat));
  OAI21_X1  g484(.A(G64gat), .B1(new_n674_), .B2(new_n368_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT48), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n368_), .A2(G64gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n680_), .B2(new_n688_), .ZN(G1333gat));
  OAI21_X1  g488(.A(G71gat), .B1(new_n674_), .B2(new_n582_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT49), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n582_), .A2(G71gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n680_), .B2(new_n692_), .ZN(G1334gat));
  OAI21_X1  g492(.A(G78gat), .B1(new_n674_), .B2(new_n375_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n375_), .A2(G78gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n680_), .B2(new_n697_), .ZN(G1335gat));
  NAND2_X1  g497(.A1(new_n679_), .A2(new_n625_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(G85gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n573_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n678_), .A2(new_n568_), .A3(new_n530_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n639_), .A2(new_n287_), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n701_), .B2(new_n705_), .ZN(G1336gat));
  NAND3_X1  g505(.A1(new_n700_), .A2(new_n355_), .A3(new_n602_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n639_), .A2(new_n368_), .A3(new_n704_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n355_), .B2(new_n708_), .ZN(G1337gat));
  NAND2_X1  g508(.A1(new_n240_), .A2(new_n414_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n639_), .A2(new_n582_), .A3(new_n704_), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n699_), .A2(new_n710_), .B1(new_n423_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g512(.A(new_n668_), .B(new_n703_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT113), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(G106gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G106gat), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n716_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT53), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n679_), .A2(new_n415_), .A3(new_n668_), .A4(new_n625_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n717_), .A2(new_n718_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .A4(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT53), .B1(new_n725_), .B2(new_n719_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1339gat));
  INV_X1    g526(.A(new_n517_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n525_), .B1(new_n519_), .B2(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT117), .ZN(new_n730_));
  AOI22_X1  g529(.A1(new_n729_), .A2(KEYINPUT117), .B1(new_n516_), .B2(new_n728_), .ZN(new_n731_));
  AOI22_X1  g530(.A1(new_n526_), .A2(new_n527_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n490_), .A2(KEYINPUT118), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n489_), .B2(new_n488_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT118), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n530_), .A2(new_n487_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n473_), .B1(new_n481_), .B2(KEYINPUT12), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n471_), .A2(KEYINPUT69), .A3(new_n464_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n740_), .A2(new_n466_), .A3(new_n741_), .A4(new_n468_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n739_), .B1(new_n742_), .B2(new_n477_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n469_), .A2(new_n475_), .A3(KEYINPUT55), .A4(new_n478_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n477_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT115), .ZN(new_n747_));
  INV_X1    g546(.A(new_n486_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n743_), .A2(new_n744_), .A3(new_n749_), .A4(new_n745_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n748_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n486_), .B1(new_n746_), .B2(KEYINPUT115), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT56), .A3(new_n750_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n738_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n737_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n738_), .ZN(new_n759_));
  AND4_X1   g558(.A1(KEYINPUT56), .A2(new_n747_), .A3(new_n748_), .A4(new_n750_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n750_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(KEYINPUT116), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n585_), .B1(new_n758_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n762_), .A2(KEYINPUT116), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n753_), .A2(new_n755_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n757_), .A3(new_n759_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n769_), .A3(new_n737_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n765_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n732_), .A2(new_n487_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n773_), .A2(KEYINPUT58), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n553_), .B1(new_n773_), .B2(KEYINPUT58), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n770_), .A2(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n568_), .B1(new_n766_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n531_), .A2(new_n568_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT114), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n678_), .A2(new_n779_), .A3(new_n553_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT54), .Z(new_n781_));
  NOR2_X1   g580(.A1(new_n777_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT59), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n573_), .B(new_n240_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n784_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n531_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n771_), .B1(new_n758_), .B2(new_n763_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n774_), .A2(new_n775_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT57), .B1(new_n770_), .B2(new_n585_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n766_), .A2(new_n776_), .A3(KEYINPUT119), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n569_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n781_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n785_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n787_), .B(new_n789_), .C1(new_n799_), .C2(new_n784_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n801_), .B(G113gat), .C1(new_n799_), .C2(new_n530_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n797_), .A2(new_n798_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n530_), .A3(new_n786_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT120), .B1(new_n804_), .B2(new_n788_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n800_), .B1(new_n802_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n800_), .B(KEYINPUT121), .C1(new_n802_), .C2(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1340gat));
  XOR2_X1   g609(.A(KEYINPUT122), .B(G120gat), .Z(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n799_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT59), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n787_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n812_), .B1(new_n815_), .B2(new_n678_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n494_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n819_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n820_), .B(new_n821_), .C1(KEYINPUT60), .C2(new_n811_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n816_), .B1(new_n813_), .B2(new_n822_), .ZN(G1341gat));
  OAI21_X1  g622(.A(G127gat), .B1(new_n815_), .B2(new_n569_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n569_), .A2(G127gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n813_), .B2(new_n825_), .ZN(G1342gat));
  INV_X1    g625(.A(G134gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n813_), .B2(new_n585_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n829_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n815_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n553_), .A2(new_n827_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n830_), .A2(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(G1343gat));
  AOI21_X1  g633(.A(new_n240_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(new_n668_), .A3(new_n368_), .A4(new_n573_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n531_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n678_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g639(.A1(new_n836_), .A2(new_n569_), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT61), .B(G155gat), .Z(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  OAI21_X1  g642(.A(G162gat), .B1(new_n836_), .B2(new_n553_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n585_), .A2(G162gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n836_), .B2(new_n845_), .ZN(G1347gat));
  NOR2_X1   g645(.A1(new_n573_), .A2(new_n368_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n240_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n668_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n782_), .A2(KEYINPUT125), .A3(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT125), .B1(new_n782_), .B2(new_n850_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n851_), .A2(new_n223_), .A3(new_n530_), .A4(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n783_), .A2(new_n530_), .A3(new_n849_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n854_), .A2(new_n855_), .A3(G169gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n854_), .B2(G169gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT126), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n853_), .B(new_n860_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1348gat));
  AND2_X1   g661(.A1(new_n851_), .A2(new_n852_), .ZN(new_n863_));
  AOI21_X1  g662(.A(G176gat), .B1(new_n863_), .B2(new_n494_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n668_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n848_), .A2(new_n678_), .A3(new_n211_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  NOR2_X1   g666(.A1(new_n848_), .A2(new_n569_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G183gat), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n569_), .A2(new_n219_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n863_), .B2(new_n870_), .ZN(G1350gat));
  NAND2_X1  g670(.A1(new_n863_), .A2(new_n554_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G190gat), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n863_), .A2(new_n548_), .A3(new_n551_), .A4(new_n215_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1351gat));
  AND4_X1   g674(.A1(new_n668_), .A2(new_n803_), .A3(new_n582_), .A4(new_n847_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(G197gat), .A3(new_n530_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT127), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n876_), .A2(new_n879_), .A3(G197gat), .A4(new_n530_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n835_), .A2(new_n668_), .A3(new_n847_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n294_), .B1(new_n881_), .B2(new_n531_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n878_), .A2(new_n880_), .A3(new_n882_), .ZN(G1352gat));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n678_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n295_), .ZN(G1353gat));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n886_));
  INV_X1    g685(.A(G211gat), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n876_), .B(new_n568_), .C1(new_n886_), .C2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n887_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1354gat));
  OAI21_X1  g689(.A(G218gat), .B1(new_n881_), .B2(new_n553_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n585_), .A2(G218gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n881_), .B2(new_n892_), .ZN(G1355gat));
endmodule


