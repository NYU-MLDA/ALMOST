//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G71gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G15gat), .B(G43gat), .Z(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT26), .B1(new_n212_), .B2(KEYINPUT82), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(G190gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n211_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n217_), .A2(new_n221_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n228_));
  INV_X1    g027(.A(new_n220_), .ZN(new_n229_));
  INV_X1    g028(.A(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n212_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT22), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(new_n223_), .A3(G169gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n222_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n227_), .A2(new_n228_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n228_), .B1(new_n227_), .B2(new_n238_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n210_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT86), .ZN(new_n244_));
  INV_X1    g043(.A(new_n218_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n226_), .A2(new_n245_), .A3(new_n229_), .A4(new_n232_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G183gat), .ZN(new_n249_));
  AND4_X1   g048(.A1(new_n247_), .A2(new_n213_), .A3(new_n216_), .A4(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n238_), .B1(new_n246_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT83), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n227_), .A2(new_n228_), .A3(new_n238_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT30), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n208_), .A2(new_n209_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n208_), .A2(new_n209_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT87), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n260_));
  INV_X1    g059(.A(G134gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G127gat), .ZN(new_n262_));
  INV_X1    g061(.A(G127gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(G134gat), .ZN(new_n264_));
  INV_X1    g063(.A(G120gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G113gat), .ZN(new_n266_));
  INV_X1    g065(.A(G113gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G120gat), .ZN(new_n268_));
  AND4_X1   g067(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .A4(new_n268_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n262_), .A2(new_n264_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n260_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n262_), .A2(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .A4(new_n268_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT88), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT31), .Z(new_n278_));
  INV_X1    g077(.A(KEYINPUT89), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n244_), .A2(new_n259_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n279_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n244_), .A2(new_n282_), .A3(new_n259_), .A4(new_n280_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n288_));
  OR2_X1    g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT90), .B1(new_n287_), .B2(KEYINPUT1), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT91), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(KEYINPUT1), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT90), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT91), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n287_), .A2(KEYINPUT1), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n289_), .A2(new_n287_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n302_), .B(KEYINPUT3), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n300_), .B(KEYINPUT2), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n277_), .B1(new_n304_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n269_), .A2(new_n270_), .ZN(new_n311_));
  AOI211_X1 g110(.A(new_n311_), .B(new_n308_), .C1(new_n299_), .C2(new_n303_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT4), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT4), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n308_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(new_n277_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G1gat), .B(G29gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G85gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT0), .B(G57gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n311_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n304_), .A2(new_n326_), .A3(new_n309_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n327_), .B(new_n318_), .C1(new_n277_), .C2(new_n315_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT101), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n310_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n331_), .A2(KEYINPUT101), .A3(new_n318_), .A4(new_n327_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n320_), .A2(new_n325_), .A3(new_n330_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n332_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n318_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n324_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n286_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n315_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT28), .B1(new_n339_), .B2(KEYINPUT29), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n339_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n342_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n343_), .B1(new_n346_), .B2(new_n340_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT92), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n344_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT92), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n339_), .A2(KEYINPUT29), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT96), .ZN(new_n354_));
  INV_X1    g153(.A(G218gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G211gat), .ZN(new_n356_));
  INV_X1    g155(.A(G211gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G218gat), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n356_), .A2(new_n358_), .A3(KEYINPUT95), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT95), .B1(new_n356_), .B2(new_n358_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n354_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT21), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT94), .B(G204gat), .ZN(new_n364_));
  AOI211_X1 g163(.A(new_n362_), .B(new_n363_), .C1(new_n364_), .C2(G197gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT95), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n357_), .A2(G218gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n355_), .A2(G211gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n356_), .A2(new_n358_), .A3(KEYINPUT95), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(KEYINPUT96), .A3(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n361_), .A2(new_n365_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n370_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n362_), .B1(G197gat), .B2(G204gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n364_), .B2(G197gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n363_), .B1(new_n364_), .B2(G197gat), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n373_), .B(new_n375_), .C1(KEYINPUT21), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n353_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT97), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n372_), .A2(new_n382_), .A3(new_n377_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n380_), .B(KEYINPUT93), .Z(new_n385_));
  NOR3_X1   g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n379_), .A2(new_n381_), .B1(new_n386_), .B2(new_n353_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n387_), .A2(new_n389_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n348_), .B(new_n352_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n387_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT98), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n388_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n345_), .A2(new_n347_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT98), .B1(new_n387_), .B2(new_n389_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n396_), .A2(new_n390_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n393_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT106), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT19), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n372_), .A2(new_n377_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n224_), .A2(new_n225_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT100), .B(KEYINPUT24), .ZN(new_n406_));
  MUX2_X1   g205(.A(new_n405_), .B(new_n224_), .S(new_n406_), .Z(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT26), .B(G190gat), .ZN(new_n408_));
  AOI211_X1 g207(.A(new_n220_), .B(new_n219_), .C1(new_n211_), .C2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n407_), .A2(new_n409_), .B1(new_n233_), .B2(new_n237_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n404_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT20), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT105), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n383_), .A2(new_n384_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n254_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n412_), .A2(new_n413_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n403_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n378_), .A2(KEYINPUT97), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n372_), .A2(new_n377_), .A3(new_n382_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n254_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT20), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT99), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n241_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT99), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT20), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n404_), .A2(new_n410_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n419_), .B1(new_n403_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT18), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n433_), .B(new_n434_), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n431_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n430_), .A2(new_n403_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n403_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n411_), .A2(KEYINPUT20), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n415_), .B2(new_n254_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n435_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n437_), .A2(KEYINPUT27), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n435_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n436_), .B(new_n441_), .C1(new_n430_), .C2(new_n403_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n401_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n444_), .A2(new_n401_), .A3(new_n448_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n338_), .B(new_n400_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n337_), .B1(new_n393_), .B2(new_n399_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n452_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n334_), .A2(new_n335_), .A3(new_n324_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT102), .B1(new_n454_), .B2(KEYINPUT33), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT102), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n333_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n446_), .A2(new_n447_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n331_), .A2(new_n319_), .A3(new_n327_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n324_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n318_), .B2(new_n317_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n463_), .B1(new_n454_), .B2(KEYINPUT33), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n459_), .A2(new_n460_), .A3(KEYINPUT103), .A4(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT103), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n425_), .A2(KEYINPUT20), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n428_), .B1(new_n467_), .B2(KEYINPUT99), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n439_), .B1(new_n468_), .B2(new_n427_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n436_), .B1(new_n469_), .B2(new_n441_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n464_), .A3(new_n443_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n455_), .A2(new_n458_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n466_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n431_), .A2(KEYINPUT32), .A3(new_n435_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n435_), .A2(KEYINPUT32), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT104), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n438_), .A2(new_n442_), .A3(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n337_), .A3(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n465_), .A2(new_n473_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n453_), .B1(new_n479_), .B2(new_n400_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n286_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n451_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G78gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(KEYINPUT68), .ZN(new_n485_));
  INV_X1    g284(.A(G64gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G57gat), .ZN(new_n487_));
  INV_X1    g286(.A(G57gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G64gat), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n487_), .A2(new_n489_), .A3(KEYINPUT68), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT11), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n483_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT11), .B1(new_n485_), .B2(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT69), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n495_), .A2(KEYINPUT69), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n495_), .A2(KEYINPUT69), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT9), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(G85gat), .A3(G92gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G85gat), .B(G92gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n503_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G106gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n511_));
  NAND2_X1  g310(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n509_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT6), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT65), .B(new_n504_), .C1(new_n505_), .C2(new_n503_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n508_), .A2(new_n515_), .A3(new_n517_), .A4(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT7), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n205_), .B(new_n509_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n522_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n517_), .A2(new_n520_), .A3(new_n523_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  INV_X1    g325(.A(new_n505_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n519_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n502_), .A2(KEYINPUT12), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(KEYINPUT67), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n533_), .B(new_n519_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n532_), .A2(new_n534_), .B1(new_n501_), .B2(new_n499_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n531_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n532_), .A2(new_n534_), .A3(new_n501_), .A4(new_n499_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G230gat), .A2(G233gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n499_), .A2(new_n501_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n545_), .A2(KEYINPUT70), .A3(new_n532_), .A4(new_n534_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT71), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n544_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n532_), .A2(new_n534_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n502_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n540_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n542_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G120gat), .B(G148gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT5), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n535_), .B1(new_n547_), .B2(KEYINPUT71), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n540_), .B1(new_n562_), .B2(new_n550_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n559_), .B1(new_n563_), .B2(new_n542_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT13), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n564_), .A3(KEYINPUT13), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G29gat), .B(G36gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G43gat), .B(G50gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT15), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573_));
  INV_X1    g372(.A(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(G8gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G1gat), .B(G8gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n571_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n579_), .B(new_n582_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(G229gat), .A3(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G113gat), .B(G141gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT80), .ZN(new_n589_));
  XOR2_X1   g388(.A(G169gat), .B(G197gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n587_), .B(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT81), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n568_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n482_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT75), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n532_), .A2(new_n571_), .A3(new_n534_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n530_), .A2(new_n572_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n601_));
  NAND2_X1  g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT74), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n598_), .A2(new_n599_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n598_), .A2(KEYINPUT74), .A3(new_n599_), .A4(new_n608_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT36), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n614_), .A2(KEYINPUT36), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n610_), .B(new_n616_), .C1(KEYINPUT36), .C2(new_n614_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT37), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n597_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n620_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(KEYINPUT75), .A3(KEYINPUT37), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(KEYINPUT76), .A3(new_n622_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT76), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n624_), .B2(KEYINPUT37), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n623_), .A2(new_n625_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G127gat), .B(G155gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT78), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n502_), .B(new_n579_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT77), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n638_), .B(new_n640_), .ZN(new_n641_));
  AOI211_X1 g440(.A(new_n637_), .B(new_n641_), .C1(new_n636_), .C2(new_n634_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n637_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n629_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n596_), .A2(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n647_), .A2(new_n574_), .A3(new_n337_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n621_), .B(KEYINPUT107), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT108), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n645_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n596_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n337_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1324gat));
  NOR2_X1   g458(.A1(new_n450_), .A2(new_n449_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n647_), .A2(new_n575_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G8gat), .B1(new_n653_), .B2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(KEYINPUT39), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(KEYINPUT39), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n666_), .B(new_n667_), .Z(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n653_), .B2(new_n286_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT41), .Z(new_n670_));
  INV_X1    g469(.A(G15gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n647_), .A2(new_n671_), .A3(new_n481_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1326gat));
  OAI21_X1  g472(.A(G22gat), .B1(new_n653_), .B2(new_n400_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT42), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n400_), .A2(G22gat), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT111), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n647_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(G1327gat));
  NOR2_X1   g478(.A1(new_n650_), .A2(new_n644_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n596_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n337_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n482_), .A2(new_n629_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n482_), .A2(new_n686_), .A3(new_n629_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n595_), .A3(new_n645_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n688_), .A2(KEYINPUT44), .A3(new_n595_), .A4(new_n645_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n337_), .A2(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n683_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n691_), .A2(new_n660_), .A3(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n681_), .A2(G36gat), .A3(new_n662_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(new_n700_), .A3(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  NAND4_X1  g504(.A1(new_n691_), .A2(G43gat), .A3(new_n481_), .A4(new_n692_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n681_), .A2(new_n286_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(G43gat), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g508(.A1(new_n681_), .A2(G50gat), .A3(new_n400_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n400_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n691_), .A2(new_n711_), .A3(new_n692_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(KEYINPUT113), .ZN(new_n713_));
  OAI21_X1  g512(.A(G50gat), .B1(new_n712_), .B2(KEYINPUT113), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(G1331gat));
  INV_X1    g514(.A(new_n568_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n593_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(new_n482_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n646_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n337_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n722_), .A2(KEYINPUT115), .A3(new_n488_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT115), .B1(new_n722_), .B2(new_n488_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n718_), .A2(new_n652_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(G57gat), .A3(new_n337_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT116), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n723_), .A2(new_n724_), .A3(new_n727_), .ZN(G1332gat));
  AOI21_X1  g527(.A(new_n486_), .B1(new_n725_), .B2(new_n660_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT48), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n721_), .A2(new_n486_), .A3(new_n660_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1333gat));
  AOI21_X1  g531(.A(new_n203_), .B1(new_n725_), .B2(new_n481_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT49), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n721_), .A2(new_n203_), .A3(new_n481_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n725_), .B2(new_n711_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT50), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n721_), .A2(new_n737_), .A3(new_n711_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1335gat));
  NOR3_X1   g540(.A1(new_n716_), .A2(new_n593_), .A3(new_n644_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT117), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(KEYINPUT117), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n654_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n718_), .A2(new_n680_), .ZN(new_n750_));
  INV_X1    g549(.A(G85gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n337_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1336gat));
  OAI21_X1  g552(.A(G92gat), .B1(new_n748_), .B2(new_n662_), .ZN(new_n754_));
  INV_X1    g553(.A(G92gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(new_n755_), .A3(new_n660_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1337gat));
  OR2_X1    g556(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n758_));
  OAI21_X1  g557(.A(G99gat), .B1(new_n748_), .B2(new_n286_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n513_), .A2(new_n514_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n286_), .A2(new_n760_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n750_), .A2(new_n761_), .B1(KEYINPUT118), .B2(KEYINPUT51), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n758_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n744_), .A2(KEYINPUT117), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n286_), .B1(new_n764_), .B2(new_n745_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n758_), .B(new_n762_), .C1(new_n765_), .C2(new_n205_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n763_), .A2(new_n767_), .ZN(G1338gat));
  AND3_X1   g567(.A1(new_n482_), .A2(new_n686_), .A3(new_n629_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n686_), .B1(new_n482_), .B2(new_n629_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n711_), .B(new_n742_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G106gat), .B1(new_n771_), .B2(KEYINPUT119), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT119), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n744_), .B2(new_n711_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT52), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n744_), .A2(new_n773_), .A3(new_n711_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n771_), .A2(KEYINPUT119), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .A4(G106gat), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n750_), .A2(new_n509_), .A3(new_n711_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n784_), .A3(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  NOR2_X1   g585(.A1(new_n660_), .A2(new_n711_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n337_), .A3(new_n481_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT123), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n591_), .B1(new_n585_), .B2(new_n581_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n580_), .A2(new_n583_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n581_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n584_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n555_), .B2(new_n560_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n554_), .B1(new_n547_), .B2(new_n538_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n541_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n552_), .A2(new_n536_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(KEYINPUT55), .A4(new_n531_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n797_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n559_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n559_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n796_), .A2(KEYINPUT121), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT121), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n563_), .A2(new_n542_), .A3(new_n559_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n795_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT58), .B1(new_n808_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n623_), .A2(new_n625_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n626_), .A2(new_n628_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n790_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n795_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n561_), .A2(KEYINPUT121), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n806_), .A2(new_n807_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n811_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(KEYINPUT122), .A3(new_n629_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n808_), .A2(KEYINPUT58), .A3(new_n811_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n816_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n807_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n559_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n561_), .B(new_n593_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n795_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  AOI211_X1 g630(.A(KEYINPUT120), .B(new_n795_), .C1(new_n561_), .C2(new_n564_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n650_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT57), .B(new_n650_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n789_), .B1(new_n825_), .B2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n816_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(KEYINPUT123), .A3(new_n835_), .A4(new_n836_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n645_), .A3(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n568_), .A2(new_n593_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n646_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT54), .ZN(new_n844_));
  AOI211_X1 g643(.A(new_n594_), .B(new_n788_), .C1(new_n841_), .C2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT124), .B1(new_n845_), .B2(G113gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n788_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n593_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n267_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n825_), .A2(new_n837_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n844_), .B1(new_n851_), .B2(new_n644_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  INV_X1    g652(.A(new_n788_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n594_), .A2(new_n267_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n855_), .B(new_n856_), .C1(new_n847_), .C2(new_n853_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n846_), .A2(new_n850_), .A3(new_n857_), .ZN(G1340gat));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n847_), .B2(new_n853_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G120gat), .B1(new_n859_), .B2(new_n716_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n265_), .B1(new_n716_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n847_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n265_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1341gat));
  OAI21_X1  g662(.A(G127gat), .B1(new_n859_), .B2(new_n645_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n847_), .A2(new_n263_), .A3(new_n644_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1342gat));
  OAI21_X1  g665(.A(G134gat), .B1(new_n859_), .B2(new_n815_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n847_), .A2(new_n261_), .A3(new_n651_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1343gat));
  AOI21_X1  g668(.A(new_n481_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n660_), .A2(new_n654_), .A3(new_n400_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n593_), .A3(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT125), .B(G141gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1344gat));
  NAND3_X1  g673(.A1(new_n870_), .A2(new_n568_), .A3(new_n871_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g675(.A1(new_n870_), .A2(new_n644_), .A3(new_n871_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  NAND2_X1  g678(.A1(new_n870_), .A2(new_n871_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G162gat), .B1(new_n880_), .B2(new_n815_), .ZN(new_n881_));
  INV_X1    g680(.A(G162gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n651_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n880_), .B2(new_n883_), .ZN(G1347gat));
  NAND2_X1  g683(.A1(new_n660_), .A2(new_n338_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n711_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n852_), .A2(new_n593_), .A3(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT62), .B1(new_n887_), .B2(KEYINPUT22), .ZN(new_n888_));
  OAI21_X1  g687(.A(G169gat), .B1(new_n887_), .B2(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n222_), .B2(new_n888_), .ZN(G1348gat));
  AND2_X1   g690(.A1(new_n852_), .A2(new_n886_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G176gat), .B1(new_n892_), .B2(new_n568_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n711_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n716_), .A2(new_n223_), .A3(new_n885_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NAND4_X1  g695(.A1(new_n894_), .A2(new_n660_), .A3(new_n338_), .A4(new_n644_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n645_), .A2(new_n211_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n897_), .A2(new_n230_), .B1(new_n892_), .B2(new_n898_), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n408_), .A3(new_n651_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n892_), .A2(new_n629_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n902_), .B2(new_n212_), .ZN(G1351gat));
  AND2_X1   g702(.A1(new_n660_), .A2(new_n452_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n870_), .A2(new_n593_), .A3(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT126), .B(G197gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1352gat));
  NAND2_X1  g706(.A1(new_n841_), .A2(new_n844_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n908_), .A2(new_n568_), .A3(new_n286_), .A4(new_n904_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G204gat), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n909_), .A2(KEYINPUT127), .A3(G204gat), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n909_), .A2(new_n364_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(G1353gat));
  XNOR2_X1  g714(.A(KEYINPUT63), .B(G211gat), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n870_), .A2(new_n644_), .A3(new_n904_), .A4(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n870_), .A2(new_n904_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n645_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n917_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  OAI21_X1  g720(.A(G218gat), .B1(new_n918_), .B2(new_n815_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n651_), .A2(new_n355_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n918_), .B2(new_n923_), .ZN(G1355gat));
endmodule


