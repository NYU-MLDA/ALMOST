//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_;
  INV_X1    g000(.A(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(G29gat), .ZN(new_n203_));
  INV_X1    g002(.A(G36gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT74), .ZN(new_n208_));
  INV_X1    g007(.A(G43gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT74), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(new_n210_), .A3(new_n206_), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n208_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n209_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n202_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n211_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G43gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n208_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(G50gat), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222_));
  INV_X1    g021(.A(G1gat), .ZN(new_n223_));
  INV_X1    g022(.A(G8gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT14), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G1gat), .B(G8gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n214_), .A2(new_n218_), .A3(KEYINPUT15), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n221_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n219_), .A2(new_n228_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n233_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n219_), .A2(new_n228_), .ZN(new_n236_));
  OAI211_X1 g035(.A(G229gat), .B(G233gat), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239_));
  INV_X1    g038(.A(G169gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G197gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT78), .ZN(new_n245_));
  INV_X1    g044(.A(new_n243_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n234_), .A2(new_n237_), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n238_), .A2(KEYINPUT78), .A3(new_n243_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT79), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(KEYINPUT79), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT84), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT86), .B(KEYINPUT2), .Z(new_n258_));
  INV_X1    g057(.A(KEYINPUT2), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n257_), .A2(new_n258_), .B1(new_n259_), .B2(new_n256_), .ZN(new_n260_));
  INV_X1    g059(.A(G141gat), .ZN(new_n261_));
  INV_X1    g060(.A(G148gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT85), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT3), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n255_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n255_), .B(KEYINPUT1), .ZN(new_n267_));
  OAI22_X1  g066(.A1(new_n267_), .A2(new_n266_), .B1(G141gat), .B2(G148gat), .ZN(new_n268_));
  OAI22_X1  g067(.A1(new_n265_), .A2(new_n266_), .B1(new_n257_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT87), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT28), .B1(new_n271_), .B2(KEYINPUT29), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n269_), .B(KEYINPUT87), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G22gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n202_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(G50gat), .A3(new_n278_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G211gat), .B(G218gat), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n286_), .A2(KEYINPUT88), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT88), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G197gat), .B(G204gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n292_), .B(KEYINPUT89), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n288_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(new_n290_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G228gat), .A2(G233gat), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n298_), .B(new_n299_), .C1(new_n273_), .C2(new_n275_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n298_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n269_), .A2(KEYINPUT29), .ZN(new_n302_));
  OAI211_X1 g101(.A(G228gat), .B(G233gat), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G78gat), .B(G106gat), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n285_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n300_), .A2(new_n303_), .A3(KEYINPUT90), .A4(new_n305_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n307_), .A2(new_n308_), .B1(new_n306_), .B2(new_n304_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n284_), .A2(new_n309_), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n304_), .A2(KEYINPUT91), .A3(new_n305_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n304_), .B1(KEYINPUT91), .B2(new_n305_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n283_), .A2(new_n281_), .A3(new_n311_), .A4(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT92), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT19), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT23), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(G183gat), .B2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT93), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT22), .B(G169gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n321_), .B(new_n323_), .C1(G176gat), .C2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT94), .ZN(new_n327_));
  NOR3_X1   g126(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n320_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI211_X1 g130(.A(new_n328_), .B(new_n329_), .C1(new_n322_), .C2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT25), .B(G183gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT26), .B(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n298_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT20), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n340_), .B1(new_n341_), .B2(G183gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n334_), .B(new_n342_), .C1(new_n333_), .C2(new_n340_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n332_), .A2(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n321_), .A2(KEYINPUT82), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n321_), .A2(KEYINPUT82), .ZN(new_n346_));
  INV_X1    g145(.A(G176gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT81), .B1(new_n240_), .B2(KEYINPUT22), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n347_), .B(new_n348_), .C1(new_n324_), .C2(KEYINPUT81), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n345_), .A2(new_n346_), .A3(new_n322_), .A4(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n298_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n318_), .B1(new_n339_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n298_), .A2(new_n351_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT20), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n318_), .A2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n354_), .B(new_n356_), .C1(new_n298_), .C2(new_n337_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT95), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n301_), .A2(new_n336_), .A3(new_n327_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n353_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369_));
  INV_X1    g168(.A(new_n367_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n353_), .A2(new_n358_), .A3(new_n361_), .A4(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n368_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n358_), .A2(new_n361_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT102), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n370_), .A4(new_n353_), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n376_));
  NAND4_X1  g175(.A1(new_n293_), .A2(new_n297_), .A3(new_n336_), .A4(new_n326_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n354_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n318_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n338_), .B(KEYINPUT20), .C1(new_n351_), .C2(new_n298_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(new_n318_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n367_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT101), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT101), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n384_), .A3(new_n367_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n371_), .A2(KEYINPUT102), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n375_), .A2(new_n383_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n372_), .B1(new_n387_), .B2(KEYINPUT27), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT0), .ZN(new_n391_));
  INV_X1    g190(.A(G57gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G127gat), .B(G134gat), .ZN(new_n395_));
  INV_X1    g194(.A(G113gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G120gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n271_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n399_), .A2(KEYINPUT99), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n401_));
  INV_X1    g200(.A(new_n398_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n273_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n271_), .A2(KEYINPUT97), .A3(new_n398_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n269_), .A2(new_n398_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(KEYINPUT4), .A4(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT98), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n399_), .A2(KEYINPUT99), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n400_), .A2(new_n406_), .A3(new_n408_), .A4(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n403_), .A2(new_n404_), .A3(new_n407_), .A4(new_n405_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n393_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n411_), .A3(new_n393_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n315_), .B1(new_n388_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n381_), .A2(KEYINPUT32), .A3(new_n370_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n373_), .A2(new_n353_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n414_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n417_), .B(new_n419_), .C1(new_n420_), .C2(new_n412_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n368_), .A2(new_n371_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n400_), .A2(new_n406_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n393_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .A4(new_n408_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n410_), .A2(KEYINPUT33), .A3(new_n411_), .A4(new_n393_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n423_), .A2(new_n424_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n421_), .A2(new_n430_), .A3(new_n314_), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n398_), .B(KEYINPUT31), .Z(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT83), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n351_), .B(KEYINPUT30), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G15gat), .B(G43gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(G71gat), .B(G99gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n437_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n438_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n416_), .A2(new_n431_), .A3(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n315_), .A2(new_n388_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n415_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n445_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n254_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT71), .ZN(new_n452_));
  NOR2_X1   g251(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n453_));
  INV_X1    g252(.A(G99gat), .ZN(new_n454_));
  INV_X1    g253(.A(G106gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  OAI22_X1  g255(.A1(KEYINPUT68), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n458_), .A2(KEYINPUT6), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(KEYINPUT6), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n456_), .B(new_n457_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  INV_X1    g261(.A(G92gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(KEYINPUT69), .A3(new_n465_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT8), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n461_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  OAI22_X1  g274(.A1(new_n475_), .A2(G106gat), .B1(new_n459_), .B2(new_n460_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n465_), .A2(KEYINPUT65), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT65), .B1(new_n465_), .B2(new_n477_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT66), .B1(G85gat), .B2(G92gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(KEYINPUT66), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT67), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  AND4_X1   g285(.A1(KEYINPUT66), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n482_), .B2(new_n481_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n465_), .A2(new_n477_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n465_), .A2(KEYINPUT65), .A3(new_n477_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n476_), .B1(new_n486_), .B2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n452_), .B(KEYINPUT12), .C1(new_n474_), .C2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G71gat), .B(G78gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(G57gat), .A2(G64gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G57gat), .A2(G64gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(KEYINPUT70), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n499_), .B1(new_n506_), .B2(KEYINPUT11), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT11), .ZN(new_n508_));
  AOI211_X1 g307(.A(new_n508_), .B(new_n498_), .C1(new_n502_), .C2(new_n505_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n486_), .A2(new_n495_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n476_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n461_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n470_), .B1(new_n461_), .B2(new_n466_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n497_), .A2(new_n512_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n518_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(new_n452_), .A3(new_n511_), .A4(KEYINPUT12), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G230gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT64), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT72), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n527_), .B1(new_n522_), .B2(new_n511_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n511_), .B2(new_n522_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n524_), .A2(KEYINPUT72), .A3(new_n527_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n530_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G176gat), .B(G204gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G120gat), .B(G148gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  AND2_X1   g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n534_), .A2(new_n539_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n451_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n511_), .B(new_n229_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT77), .Z(new_n550_));
  XNOR2_X1  g349(.A(G127gat), .B(G155gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT16), .ZN(new_n552_));
  INV_X1    g351(.A(G183gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT17), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n549_), .A2(new_n452_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n549_), .A2(new_n452_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n221_), .A2(new_n522_), .A3(new_n230_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n219_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT34), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT35), .Z(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT75), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n568_), .A2(new_n569_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(KEYINPUT35), .A3(new_n571_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n574_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n567_), .B1(new_n579_), .B2(KEYINPUT36), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n567_), .A2(KEYINPUT36), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n583_), .B(new_n579_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(KEYINPUT37), .A3(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n546_), .A2(new_n563_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n223_), .A3(new_n415_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n587_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n563_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n545_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n250_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n597_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n223_), .B1(new_n601_), .B2(new_n415_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n595_), .A2(new_n602_), .ZN(G1324gat));
  NAND3_X1  g402(.A1(new_n592_), .A2(new_n224_), .A3(new_n388_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n388_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G8gat), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n606_), .A2(KEYINPUT39), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(KEYINPUT39), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g409(.A(G15gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n601_), .B2(new_n449_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT41), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n592_), .A2(new_n611_), .A3(new_n449_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1326gat));
  NAND3_X1  g414(.A1(new_n592_), .A2(new_n277_), .A3(new_n315_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n277_), .B1(new_n601_), .B2(new_n315_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n619_), .A2(KEYINPUT42), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT42), .B1(new_n619_), .B2(new_n620_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n616_), .B1(new_n621_), .B2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n591_), .ZN(new_n624_));
  AOI211_X1 g423(.A(KEYINPUT43), .B(new_n624_), .C1(new_n446_), .C2(new_n450_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT43), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n446_), .A2(new_n450_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n627_), .B2(new_n591_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n563_), .B(new_n600_), .C1(new_n625_), .C2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT44), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n591_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT43), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n627_), .A2(new_n626_), .A3(new_n591_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n635_), .A2(KEYINPUT44), .A3(new_n563_), .A4(new_n600_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G29gat), .B1(new_n637_), .B2(new_n448_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n546_), .A2(new_n598_), .A3(new_n587_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n203_), .A3(new_n415_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1328gat));
  NAND3_X1  g440(.A1(new_n631_), .A2(new_n636_), .A3(new_n388_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n587_), .A2(new_n598_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n451_), .A2(new_n204_), .A3(new_n545_), .A4(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n388_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n646_));
  OR3_X1    g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n648_));
  AOI22_X1  g447(.A1(new_n642_), .A2(G36gat), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT106), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT106), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n649_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  NAND3_X1  g454(.A1(new_n631_), .A2(new_n636_), .A3(new_n449_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G43gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n639_), .A2(new_n209_), .A3(new_n449_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT47), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1330gat));
  OAI21_X1  g460(.A(G50gat), .B1(new_n637_), .B2(new_n314_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n639_), .A2(new_n202_), .A3(new_n315_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1331gat));
  NOR2_X1   g463(.A1(new_n545_), .A2(new_n251_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n627_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n591_), .A2(new_n563_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n415_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n563_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n597_), .A2(new_n599_), .A3(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT107), .Z(new_n673_));
  NOR2_X1   g472(.A1(new_n448_), .A2(new_n392_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(G1332gat));
  OR3_X1    g474(.A1(new_n668_), .A2(G64gat), .A3(new_n645_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n388_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT48), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n677_), .A2(new_n678_), .A3(G64gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n677_), .B2(G64gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(G1333gat));
  OR3_X1    g480(.A1(new_n668_), .A2(G71gat), .A3(new_n445_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n673_), .A2(new_n449_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G71gat), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT49), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT49), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1334gat));
  NAND2_X1  g486(.A1(new_n673_), .A2(new_n315_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G78gat), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(KEYINPUT50), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(KEYINPUT50), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n314_), .A2(G78gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT108), .ZN(new_n693_));
  OAI22_X1  g492(.A1(new_n690_), .A2(new_n691_), .B1(new_n668_), .B2(new_n693_), .ZN(G1335gat));
  NAND2_X1  g493(.A1(new_n666_), .A2(new_n643_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT109), .Z(new_n696_));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n415_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n665_), .A2(new_n563_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT110), .Z(new_n699_));
  AND2_X1   g498(.A1(new_n635_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n448_), .A2(new_n462_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1336gat));
  AOI21_X1  g501(.A(G92gat), .B1(new_n696_), .B2(new_n388_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n645_), .A2(new_n463_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n700_), .B2(new_n704_), .ZN(G1337gat));
  AOI21_X1  g504(.A(new_n454_), .B1(new_n700_), .B2(new_n449_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n445_), .A2(new_n475_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n696_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT51), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(G1338gat));
  OAI211_X1 g509(.A(new_n699_), .B(new_n315_), .C1(new_n625_), .C2(new_n628_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G106gat), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT111), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n714_), .A3(G106gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(KEYINPUT52), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n696_), .A2(new_n455_), .A3(new_n315_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n712_), .A2(KEYINPUT111), .A3(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT53), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT53), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n716_), .A2(new_n717_), .A3(new_n722_), .A4(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1339gat));
  INV_X1    g523(.A(KEYINPUT116), .ZN(new_n725_));
  INV_X1    g524(.A(new_n447_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n250_), .A2(new_n541_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  INV_X1    g527(.A(new_n539_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n526_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n529_), .B1(KEYINPUT112), .B2(KEYINPUT55), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n730_), .B2(KEYINPUT72), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n734_), .B2(KEYINPUT55), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n524_), .A2(new_n527_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n728_), .B(new_n729_), .C1(new_n735_), .C2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT55), .B1(new_n533_), .B2(KEYINPUT112), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n730_), .A2(new_n731_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT56), .B1(new_n741_), .B2(new_n539_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n727_), .B1(new_n738_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT113), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n232_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n231_), .A2(new_n233_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n745_), .B(new_n243_), .C1(new_n746_), .C2(new_n232_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n247_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n529_), .B(new_n526_), .C1(new_n521_), .C2(new_n523_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n733_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n736_), .B1(new_n752_), .B2(new_n732_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n728_), .B1(new_n753_), .B2(new_n729_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n741_), .A2(KEYINPUT56), .A3(new_n539_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n727_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n744_), .A2(new_n749_), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT57), .A3(new_n587_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT115), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n587_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n541_), .B1(new_n742_), .B2(KEYINPUT114), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n765_), .A2(KEYINPUT58), .A3(new_n748_), .A4(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n766_), .B(new_n748_), .C1(KEYINPUT114), .C2(new_n756_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n591_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n759_), .A2(new_n772_), .A3(KEYINPUT57), .A4(new_n587_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n761_), .A2(new_n764_), .A3(new_n771_), .A4(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n563_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n589_), .A2(new_n545_), .A3(new_n671_), .A4(new_n590_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n726_), .B1(new_n775_), .B2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n448_), .A2(new_n445_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n725_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n778_), .B1(new_n774_), .B2(new_n563_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n781_), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n783_), .A2(KEYINPUT116), .A3(new_n726_), .A4(new_n784_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G113gat), .B1(new_n786_), .B2(new_n251_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n789_));
  NOR4_X1   g588(.A1(new_n783_), .A2(KEYINPUT59), .A3(new_n726_), .A4(new_n784_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n254_), .A2(new_n396_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n787_), .B1(new_n791_), .B2(new_n792_), .ZN(G1340gat));
  INV_X1    g592(.A(G120gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT60), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n545_), .B2(G120gat), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n795_), .B(new_n797_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n789_), .A2(new_n790_), .A3(new_n545_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n794_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT117), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n798_), .B(new_n802_), .C1(new_n799_), .C2(new_n794_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1341gat));
  AOI21_X1  g603(.A(G127gat), .B1(new_n786_), .B2(new_n598_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n598_), .A2(G127gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n791_), .B2(new_n806_), .ZN(G1342gat));
  AOI21_X1  g606(.A(G134gat), .B1(new_n786_), .B2(new_n596_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n591_), .A2(G134gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n791_), .B2(new_n809_), .ZN(G1343gat));
  NOR2_X1   g609(.A1(new_n449_), .A2(new_n314_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n783_), .A2(new_n448_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n645_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n250_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(new_n261_), .ZN(G1344gat));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n545_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(new_n262_), .ZN(G1345gat));
  NOR2_X1   g617(.A1(new_n814_), .A2(new_n563_), .ZN(new_n819_));
  XOR2_X1   g618(.A(KEYINPUT61), .B(G155gat), .Z(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1346gat));
  INV_X1    g620(.A(new_n814_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n822_), .A2(G162gat), .A3(new_n591_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G162gat), .B1(new_n822_), .B2(new_n596_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1347gat));
  NOR2_X1   g624(.A1(new_n783_), .A2(new_n315_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n449_), .A2(new_n448_), .A3(new_n388_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT118), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n251_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G169gat), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n834_), .B(new_n835_), .C1(new_n325_), .C2(new_n831_), .ZN(G1348gat));
  AOI21_X1  g635(.A(G176gat), .B1(new_n830_), .B2(new_n599_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n826_), .B(KEYINPUT119), .Z(new_n838_));
  AND2_X1   g637(.A1(new_n838_), .A2(new_n828_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n545_), .A2(new_n347_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(G1349gat));
  NOR3_X1   g640(.A1(new_n829_), .A2(new_n563_), .A3(new_n333_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n598_), .A3(new_n828_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n553_), .ZN(G1350gat));
  NAND2_X1  g643(.A1(new_n775_), .A2(new_n779_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n845_), .A2(new_n314_), .A3(new_n591_), .A4(new_n828_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n846_), .A2(KEYINPUT120), .A3(G190gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT120), .B1(new_n846_), .B2(G190gat), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n596_), .A2(new_n334_), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT121), .Z(new_n850_));
  OAI22_X1  g649(.A1(new_n847_), .A2(new_n848_), .B1(new_n829_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI221_X1 g652(.A(KEYINPUT122), .B1(new_n829_), .B2(new_n850_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1351gat));
  NOR2_X1   g654(.A1(new_n645_), .A2(new_n415_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n845_), .A2(new_n811_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT123), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n783_), .A2(new_n812_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n856_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n250_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT125), .B1(new_n862_), .B2(G197gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n859_), .B2(new_n856_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n856_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n783_), .A2(KEYINPUT123), .A3(new_n812_), .A4(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n251_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n242_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n862_), .A2(new_n870_), .A3(G197gat), .ZN(new_n871_));
  OAI211_X1 g670(.A(G197gat), .B(new_n251_), .C1(new_n864_), .C2(new_n866_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT124), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n863_), .A2(new_n869_), .B1(new_n871_), .B2(new_n873_), .ZN(G1352gat));
  NAND2_X1  g673(.A1(new_n858_), .A2(new_n861_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n599_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n598_), .A3(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT126), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n879_), .B(new_n881_), .ZN(G1354gat));
  NOR2_X1   g681(.A1(new_n587_), .A2(G218gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n624_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n885_));
  INV_X1    g684(.A(G218gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT127), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT127), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(new_n884_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1355gat));
endmodule


