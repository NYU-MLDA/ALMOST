//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n941_,
    new_n943_, new_n944_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G227gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(G15gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT87), .B(G43gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G71gat), .B(G99gat), .Z(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT80), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT83), .B(KEYINPUT23), .Z(new_n221_));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI22_X1  g022(.A1(new_n223_), .A2(KEYINPUT84), .B1(KEYINPUT23), .B2(new_n222_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n225_));
  INV_X1    g024(.A(new_n222_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT84), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n220_), .B1(new_n224_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT85), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n222_), .A2(KEYINPUT23), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n228_), .B2(new_n227_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT85), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n220_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n219_), .B1(G169gat), .B2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n218_), .A2(new_n238_), .A3(KEYINPUT81), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT81), .B1(new_n218_), .B2(new_n238_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT25), .B(G183gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT26), .B(G190gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT82), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n239_), .A2(new_n246_), .A3(new_n240_), .A4(new_n243_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n231_), .A2(new_n236_), .A3(new_n245_), .A4(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT86), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n249_), .B1(new_n222_), .B2(KEYINPUT23), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n225_), .A2(new_n249_), .A3(new_n226_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G169gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n248_), .A2(KEYINPUT30), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT30), .B1(new_n248_), .B2(new_n258_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT88), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n248_), .A2(new_n258_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT30), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT88), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n259_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n213_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n265_), .B2(new_n259_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n213_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n207_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n260_), .A2(new_n261_), .A3(KEYINPUT88), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(new_n273_), .B2(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n262_), .A2(new_n213_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n206_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G197gat), .B(G204gat), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT96), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G197gat), .B(G204gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT96), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G211gat), .B(G218gat), .Z(new_n284_));
  NAND4_X1  g083(.A1(new_n280_), .A2(KEYINPUT21), .A3(new_n283_), .A4(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT97), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n284_), .A2(KEYINPUT21), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n288_), .A2(KEYINPUT97), .A3(new_n283_), .A4(new_n280_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n281_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n284_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n281_), .A2(KEYINPUT94), .A3(new_n291_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT94), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n279_), .B2(KEYINPUT21), .ZN(new_n297_));
  OAI221_X1 g096(.A(new_n294_), .B1(new_n293_), .B2(new_n292_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(G228gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT92), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(KEYINPUT92), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT93), .Z(new_n305_));
  AND2_X1   g104(.A1(new_n299_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G141gat), .B(G148gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n311_), .B2(KEYINPUT1), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n312_), .B2(KEYINPUT90), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT90), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n314_), .B(new_n309_), .C1(new_n311_), .C2(KEYINPUT1), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n308_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT3), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT2), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n311_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n322_), .A2(new_n309_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n316_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n307_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n323_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n313_), .A2(new_n315_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(new_n308_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n306_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n299_), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n336_));
  NOR2_X1   g135(.A1(new_n324_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n304_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n332_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT99), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n324_), .A2(new_n325_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT28), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n341_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n299_), .A2(new_n305_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n304_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n324_), .A2(new_n336_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(new_n299_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n347_), .A2(new_n333_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n334_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT100), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT100), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n333_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n339_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n345_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT100), .B1(new_n351_), .B2(new_n352_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n354_), .A3(new_n339_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n358_), .A2(new_n340_), .A3(new_n344_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n278_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT18), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  AND2_X1   g165(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT19), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n234_), .A2(new_n253_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n257_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n214_), .A2(new_n219_), .ZN(new_n373_));
  AND4_X1   g172(.A1(new_n251_), .A2(new_n254_), .A3(new_n243_), .A4(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n237_), .A2(KEYINPUT101), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n237_), .A2(KEYINPUT101), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n375_), .A2(new_n217_), .A3(new_n215_), .A4(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n299_), .B1(new_n379_), .B2(KEYINPUT105), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(KEYINPUT105), .B2(new_n379_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n263_), .B2(new_n299_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n370_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n379_), .B2(new_n299_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n263_), .B2(new_n299_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(new_n369_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n367_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n204_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n329_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT4), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OR3_X1    g192(.A1(new_n324_), .A2(new_n389_), .A3(KEYINPUT4), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT103), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT103), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n390_), .A2(new_n398_), .A3(new_n392_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n395_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G85gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G57gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n395_), .A2(new_n397_), .A3(new_n404_), .A4(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n263_), .A2(new_n299_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n371_), .A2(new_n257_), .B1(new_n377_), .B2(new_n374_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n369_), .B1(new_n335_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(KEYINPUT20), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT102), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT102), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n383_), .A2(new_n414_), .A3(new_n411_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n386_), .A2(new_n369_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n388_), .B(new_n408_), .C1(new_n417_), .C2(new_n367_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n407_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n404_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n421_), .A2(KEYINPUT104), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n391_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(KEYINPUT104), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n407_), .A2(new_n419_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n366_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n417_), .A2(new_n429_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n412_), .A2(KEYINPUT102), .B1(new_n386_), .B2(new_n369_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n366_), .A3(new_n415_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n418_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n362_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n429_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(KEYINPUT27), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT27), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT106), .B1(new_n433_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT106), .ZN(new_n440_));
  AOI211_X1 g239(.A(new_n440_), .B(KEYINPUT27), .C1(new_n430_), .C2(new_n432_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n437_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n408_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n277_), .A2(new_n361_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n276_), .A2(new_n272_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n435_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n449_));
  OR2_X1    g248(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n450_));
  INV_X1    g249(.A(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT6), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(G99gat), .A3(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT9), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(KEYINPUT64), .ZN(new_n460_));
  AND2_X1   g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n453_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G85gat), .A2(G92gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT9), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT64), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(new_n459_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n449_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n455_), .A2(new_n457_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n471_));
  AND4_X1   g270(.A1(new_n449_), .A2(new_n469_), .A3(new_n471_), .A4(new_n453_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n461_), .A2(new_n464_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n458_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n476_));
  INV_X1    g275(.A(G99gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n451_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n479_));
  OR2_X1    g278(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n474_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT67), .B(new_n474_), .C1(new_n475_), .C2(new_n481_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(KEYINPUT8), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT8), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n473_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(G71gat), .ZN(new_n491_));
  INV_X1    g290(.A(G71gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(KEYINPUT68), .ZN(new_n493_));
  OAI21_X1  g292(.A(G78gat), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(KEYINPUT68), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(G71gat), .ZN(new_n496_));
  INV_X1    g295(.A(G78gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G64gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G57gat), .ZN(new_n500_));
  INV_X1    g299(.A(G57gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G64gat), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n500_), .A2(new_n502_), .A3(KEYINPUT11), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT11), .B1(new_n500_), .B2(new_n502_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n494_), .B(new_n498_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT69), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n500_), .A2(new_n502_), .A3(KEYINPUT11), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n497_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n505_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n506_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI211_X1 g312(.A(new_n448_), .B(KEYINPUT12), .C1(new_n489_), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n485_), .A2(KEYINPUT8), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n458_), .A2(new_n479_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT67), .B1(new_n516_), .B2(new_n474_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n469_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n453_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT65), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n463_), .A2(new_n449_), .A3(new_n469_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n488_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n513_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT12), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT71), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n514_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G230gat), .A2(G233gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(new_n523_), .B2(new_n518_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n473_), .A2(new_n486_), .A3(KEYINPUT70), .A4(new_n488_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n505_), .A2(new_n510_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(new_n525_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n530_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n523_), .A2(new_n518_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(KEYINPUT69), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n505_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n527_), .A2(new_n528_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n524_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n528_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G120gat), .B(G148gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT5), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n542_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT13), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT13), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G1gat), .B(G8gat), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT76), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(G15gat), .ZN(new_n562_));
  INV_X1    g361(.A(G22gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G15gat), .A2(G22gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G1gat), .A2(G8gat), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n564_), .A2(new_n565_), .B1(KEYINPUT14), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n561_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G29gat), .B(G36gat), .Z(new_n569_));
  XOR2_X1   g368(.A(G43gat), .B(G50gat), .Z(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n561_), .A2(new_n567_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n561_), .A2(new_n567_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n571_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT77), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT77), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n579_), .A3(new_n576_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n578_), .A2(G229gat), .A3(G233gat), .A4(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n572_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT78), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n581_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G169gat), .B(G197gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT79), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT79), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n581_), .A2(new_n588_), .A3(new_n595_), .A4(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n593_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n558_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n568_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(new_n532_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  XOR2_X1   g405(.A(G127gat), .B(G155gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT16), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n605_), .A2(new_n606_), .A3(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n533_), .B2(new_n603_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n610_), .B(new_n606_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n604_), .B2(new_n539_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n614_), .B1(new_n539_), .B2(new_n604_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(KEYINPUT36), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT34), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT35), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT74), .B1(new_n623_), .B2(new_n624_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT73), .B1(new_n489_), .B2(new_n571_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT73), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n536_), .A2(new_n630_), .A3(new_n572_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n585_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n572_), .A2(new_n584_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n530_), .B(new_n531_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n626_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n632_), .A2(new_n626_), .A3(new_n635_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n620_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n620_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n636_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT36), .ZN(new_n643_));
  INV_X1    g442(.A(new_n619_), .ZN(new_n644_));
  OAI22_X1  g443(.A1(new_n639_), .A2(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT37), .B1(new_n642_), .B2(KEYINPUT75), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n641_), .B1(new_n640_), .B2(new_n636_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n637_), .A2(new_n620_), .A3(new_n638_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n648_), .A2(new_n649_), .B1(KEYINPUT36), .B2(new_n619_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT75), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n616_), .B1(new_n647_), .B2(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n447_), .A2(new_n601_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(G1gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n408_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT107), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n447_), .A2(new_n601_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n645_), .A2(new_n616_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(new_n408_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n661_), .B(new_n662_), .C1(new_n657_), .C2(new_n666_), .ZN(G1324gat));
  NAND4_X1  g466(.A1(new_n447_), .A2(new_n601_), .A3(new_n442_), .A4(new_n664_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT108), .B1(new_n668_), .B2(G8gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(KEYINPUT109), .B2(KEYINPUT39), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(KEYINPUT108), .A3(G8gat), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(new_n671_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n671_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n672_), .B(new_n673_), .C1(new_n676_), .C2(new_n669_), .ZN(new_n677_));
  INV_X1    g476(.A(G8gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n656_), .A2(new_n678_), .A3(new_n442_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n675_), .A2(new_n677_), .A3(new_n679_), .A4(new_n681_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1325gat));
  AOI21_X1  g484(.A(new_n562_), .B1(new_n665_), .B2(new_n278_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n656_), .A2(new_n562_), .A3(new_n278_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1326gat));
  AOI21_X1  g489(.A(new_n563_), .B1(new_n665_), .B2(new_n361_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT42), .Z(new_n692_));
  NAND2_X1  g491(.A1(new_n361_), .A2(new_n563_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT112), .Z(new_n694_));
  NAND2_X1  g493(.A1(new_n656_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1327gat));
  INV_X1    g495(.A(new_n616_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n650_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n663_), .A2(new_n698_), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n699_), .A2(G29gat), .A3(new_n443_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n437_), .ZN(new_n701_));
  AND4_X1   g500(.A1(new_n366_), .A2(new_n413_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n366_), .B1(new_n431_), .B2(new_n415_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n438_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n440_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n433_), .A2(KEYINPUT106), .A3(new_n438_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n277_), .A2(new_n361_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n272_), .A2(new_n357_), .A3(new_n276_), .A4(new_n360_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n408_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n707_), .A2(new_n710_), .B1(new_n434_), .B2(new_n362_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n647_), .A2(new_n654_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  INV_X1    g513(.A(new_n712_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n447_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n601_), .A2(new_n616_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n721_), .B(new_n718_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n408_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G29gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n723_), .B2(new_n408_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n700_), .B1(new_n726_), .B2(new_n727_), .ZN(G1328gat));
  OR2_X1    g527(.A1(new_n442_), .A2(KEYINPUT114), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n442_), .A2(KEYINPUT114), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n699_), .A2(new_n733_), .A3(KEYINPUT45), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT45), .B1(new_n699_), .B2(new_n733_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n720_), .A2(new_n722_), .A3(new_n707_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n732_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT115), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT116), .Z(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n741_), .B(new_n736_), .C1(new_n737_), .C2(new_n732_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  INV_X1    g544(.A(G43gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n277_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n723_), .A2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n699_), .B2(new_n277_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(KEYINPUT47), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n748_), .B2(new_n749_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1330gat));
  INV_X1    g551(.A(new_n361_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n699_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(G50gat), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n361_), .A2(G50gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n723_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1331gat));
  INV_X1    g558(.A(new_n558_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n599_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n447_), .A2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n664_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G57gat), .B1(new_n764_), .B2(new_n443_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n762_), .A2(new_n655_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n501_), .A3(new_n408_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1332gat));
  AOI21_X1  g567(.A(new_n499_), .B1(new_n763_), .B2(new_n731_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT48), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n766_), .A2(new_n499_), .A3(new_n731_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1333gat));
  AOI21_X1  g571(.A(new_n492_), .B1(new_n763_), .B2(new_n278_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT49), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n766_), .A2(new_n492_), .A3(new_n278_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1334gat));
  AOI21_X1  g575(.A(new_n497_), .B1(new_n763_), .B2(new_n361_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT50), .Z(new_n778_));
  NAND2_X1  g577(.A1(new_n361_), .A2(new_n497_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT118), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n766_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(G1335gat));
  AND2_X1   g581(.A1(new_n762_), .A2(new_n698_), .ZN(new_n783_));
  INV_X1    g582(.A(G85gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n784_), .A3(new_n408_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n761_), .A2(new_n616_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n713_), .B2(new_n716_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n408_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n785_), .B1(new_n788_), .B2(new_n784_), .ZN(G1336gat));
  INV_X1    g588(.A(G92gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n783_), .A2(new_n790_), .A3(new_n442_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n787_), .A2(new_n731_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n790_), .ZN(G1337gat));
  NAND2_X1  g592(.A1(new_n450_), .A2(new_n452_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n783_), .A2(new_n795_), .A3(new_n278_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n783_), .A2(KEYINPUT119), .A3(new_n795_), .A4(new_n278_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n787_), .A2(new_n278_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n477_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT51), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n799_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n804_), .B(new_n805_), .C1(new_n477_), .C2(new_n801_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(G1338gat));
  XNOR2_X1  g606(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n786_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n711_), .A2(KEYINPUT43), .A3(new_n712_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n714_), .B1(new_n447_), .B2(new_n715_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n361_), .B(new_n810_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(G106gat), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT52), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n813_), .B2(G106gat), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n753_), .B(new_n786_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT120), .B(new_n819_), .C1(new_n820_), .C2(new_n451_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n783_), .A2(new_n451_), .A3(new_n361_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n809_), .B1(new_n818_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT120), .B1(new_n820_), .B2(new_n451_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT52), .A3(new_n815_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(new_n821_), .A3(new_n822_), .A4(new_n808_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(G1339gat));
  AND3_X1   g627(.A1(new_n555_), .A2(new_n600_), .A3(new_n557_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n655_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n655_), .B2(new_n829_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n599_), .A2(new_n551_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n488_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n539_), .B1(new_n486_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n448_), .B1(new_n838_), .B2(KEYINPUT12), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n524_), .A2(KEYINPUT71), .A3(new_n525_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n839_), .A2(new_n540_), .A3(new_n535_), .A4(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n836_), .B1(new_n841_), .B2(new_n544_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n544_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n527_), .A2(KEYINPUT55), .A3(new_n541_), .A4(new_n528_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n549_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n528_), .B1(new_n527_), .B2(new_n541_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n542_), .B1(new_n850_), .B2(new_n836_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n845_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT56), .A3(new_n549_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n835_), .B1(new_n849_), .B2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n578_), .A2(new_n580_), .A3(new_n587_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n583_), .A2(new_n585_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n855_), .B(new_n593_), .C1(new_n856_), .C2(new_n587_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n597_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n554_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n650_), .B1(new_n854_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n858_), .A2(new_n552_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT56), .B1(new_n852_), .B2(new_n549_), .ZN(new_n864_));
  AOI211_X1 g663(.A(new_n848_), .B(new_n550_), .C1(new_n851_), .C2(new_n845_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT58), .B(new_n863_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n715_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n552_), .B1(new_n598_), .B2(new_n597_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n859_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(KEYINPUT57), .A3(new_n650_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n862_), .A2(new_n870_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n834_), .B1(new_n876_), .B2(new_n616_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n443_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n442_), .A2(new_n709_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(G113gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n599_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n880_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n878_), .A2(KEYINPUT59), .A3(new_n879_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n600_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n883_), .B1(new_n887_), .B2(new_n882_), .ZN(G1340gat));
  INV_X1    g687(.A(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n760_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n881_), .B(new_n890_), .C1(KEYINPUT60), .C2(new_n889_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n760_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g692(.A(G127gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n616_), .A2(new_n894_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n878_), .A2(KEYINPUT59), .A3(new_n879_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT59), .B1(new_n878_), .B2(new_n879_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(KEYINPUT123), .B(new_n894_), .C1(new_n880_), .C2(new_n616_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n876_), .A2(new_n616_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n834_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  AND4_X1   g702(.A1(new_n408_), .A2(new_n903_), .A3(new_n697_), .A4(new_n879_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n900_), .B1(new_n904_), .B2(G127gat), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n898_), .A2(new_n899_), .A3(new_n905_), .ZN(G1342gat));
  INV_X1    g705(.A(G134gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n881_), .A2(new_n907_), .A3(new_n645_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n712_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1343gat));
  NOR2_X1   g709(.A1(new_n731_), .A2(new_n708_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n878_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n599_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n558_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g715(.A1(new_n903_), .A2(new_n408_), .A3(new_n697_), .A4(new_n911_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT124), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n878_), .A2(new_n919_), .A3(new_n697_), .A4(new_n911_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT61), .B(G155gat), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n918_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n918_), .B2(new_n920_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1346gat));
  AOI21_X1  g723(.A(G162gat), .B1(new_n912_), .B2(new_n645_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n715_), .A2(G162gat), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT125), .Z(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n912_), .B2(new_n927_), .ZN(G1347gat));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n731_), .A2(new_n443_), .ZN(new_n930_));
  NOR4_X1   g729(.A1(new_n877_), .A2(new_n600_), .A3(new_n930_), .A4(new_n709_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT22), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n929_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G169gat), .ZN(new_n934_));
  INV_X1    g733(.A(G169gat), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n931_), .B2(new_n929_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n934_), .B1(new_n933_), .B2(new_n936_), .ZN(G1348gat));
  NOR3_X1   g736(.A1(new_n877_), .A2(new_n709_), .A3(new_n930_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n558_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n697_), .ZN(new_n941_));
  MUX2_X1   g740(.A(new_n241_), .B(G183gat), .S(new_n941_), .Z(G1350gat));
  NAND3_X1  g741(.A1(new_n938_), .A2(new_n242_), .A3(new_n645_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n938_), .A2(new_n715_), .ZN(new_n944_));
  INV_X1    g743(.A(G190gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n944_), .B2(new_n945_), .ZN(G1351gat));
  INV_X1    g745(.A(new_n930_), .ZN(new_n947_));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n874_), .B2(new_n650_), .ZN(new_n948_));
  AOI211_X1 g747(.A(new_n861_), .B(new_n645_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n697_), .B1(new_n950_), .B2(new_n870_), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n445_), .B(new_n947_), .C1(new_n951_), .C2(new_n834_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(KEYINPUT126), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n930_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n954_), .A2(new_n955_), .A3(new_n445_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n953_), .A2(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(G197gat), .B1(new_n957_), .B2(new_n599_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n955_), .B1(new_n954_), .B2(new_n445_), .ZN(new_n959_));
  NOR4_X1   g758(.A1(new_n877_), .A2(KEYINPUT126), .A3(new_n930_), .A4(new_n708_), .ZN(new_n960_));
  OAI211_X1 g759(.A(G197gat), .B(new_n599_), .C1(new_n959_), .C2(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n958_), .A2(new_n962_), .ZN(G1352gat));
  OAI21_X1  g762(.A(new_n558_), .B1(new_n959_), .B2(new_n960_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n964_), .A2(KEYINPUT127), .A3(G204gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n957_), .A2(new_n558_), .A3(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n967_), .ZN(G1353gat));
  OR2_X1    g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n969_), .B1(new_n957_), .B2(new_n697_), .ZN(new_n970_));
  XOR2_X1   g769(.A(KEYINPUT63), .B(G211gat), .Z(new_n971_));
  OAI211_X1 g770(.A(new_n697_), .B(new_n971_), .C1(new_n959_), .C2(new_n960_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n972_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n970_), .A2(new_n973_), .ZN(G1354gat));
  INV_X1    g773(.A(G218gat), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n957_), .A2(new_n975_), .A3(new_n645_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n712_), .B1(new_n953_), .B2(new_n956_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n975_), .B2(new_n977_), .ZN(G1355gat));
endmodule


