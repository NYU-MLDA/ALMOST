//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT6), .Z(new_n208_));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209_));
  AND2_X1   g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G85gat), .B(G92gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT10), .B(G99gat), .ZN(new_n213_));
  OAI221_X1 g012(.A(new_n211_), .B1(new_n209_), .B2(new_n212_), .C1(G106gat), .C2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n212_), .B(KEYINPUT64), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT7), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n217_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n208_), .A2(KEYINPUT65), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n220_), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n216_), .B1(new_n225_), .B2(new_n215_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n214_), .B1(new_n221_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n228_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G57gat), .B(G64gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT11), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT67), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(KEYINPUT11), .B2(new_n232_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT68), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n231_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n239_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(new_n227_), .A3(KEYINPUT12), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n231_), .A2(new_n240_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n241_), .B(new_n243_), .C1(new_n244_), .C2(KEYINPUT12), .ZN(new_n245_));
  AND2_X1   g044(.A1(G230gat), .A2(G233gat), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(KEYINPUT69), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n241_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n244_), .A2(KEYINPUT69), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n246_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n206_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n247_), .A2(new_n251_), .A3(new_n206_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT13), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(KEYINPUT13), .A3(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT70), .Z(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT74), .B(G1gat), .Z(new_n261_));
  INV_X1    g060(.A(G8gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT14), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G15gat), .B(G22gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G1gat), .B(G8gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT75), .Z(new_n268_));
  AND2_X1   g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n270_), .A2(new_n242_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT17), .ZN(new_n272_));
  XOR2_X1   g071(.A(G127gat), .B(G155gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT16), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G183gat), .B(G211gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n271_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n242_), .B2(new_n270_), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n270_), .B(new_n240_), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n276_), .B(new_n272_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT76), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G29gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G43gat), .B(G50gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n229_), .A2(new_n286_), .A3(new_n230_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n286_), .B(KEYINPUT15), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n227_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G232gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n287_), .A2(new_n288_), .A3(new_n290_), .A4(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n287_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n293_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT35), .B1(new_n287_), .B2(new_n290_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT72), .B(new_n295_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G190gat), .B(G218gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G134gat), .B(G162gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n299_), .B1(KEYINPUT36), .B2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n287_), .A2(new_n290_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n296_), .B(new_n293_), .C1(new_n304_), .C2(KEYINPUT35), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n302_), .A2(KEYINPUT36), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n305_), .A2(KEYINPUT72), .A3(new_n295_), .A4(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n295_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n302_), .A2(KEYINPUT36), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT37), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT37), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n303_), .A2(new_n307_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n315_), .B1(new_n316_), .B2(KEYINPUT73), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n283_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n260_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(G15gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(G71gat), .B(G99gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT82), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n328_), .B2(KEYINPUT23), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(G183gat), .B2(G190gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G169gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n334_), .B1(G183gat), .B2(G190gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n328_), .B2(new_n334_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(KEYINPUT24), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(KEYINPUT24), .A3(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT81), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n333_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n349_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n325_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n354_), .A2(new_n324_), .A3(new_n350_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n323_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n324_), .B1(new_n354_), .B2(new_n350_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n351_), .A2(new_n325_), .A3(new_n352_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n323_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT83), .B(G43gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n362_), .A3(new_n360_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT31), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT31), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n364_), .A2(new_n365_), .A3(new_n369_), .A4(new_n366_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G113gat), .B(G120gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n371_), .B(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT1), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT86), .Z(new_n379_));
  NOR2_X1   g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n377_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT89), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n381_), .A2(new_n380_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n396_));
  NOR4_X1   g195(.A1(new_n396_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT87), .B1(new_n388_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n395_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT88), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n404_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n392_), .B(new_n393_), .C1(new_n400_), .C2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n409_));
  INV_X1    g208(.A(G141gat), .ZN(new_n410_));
  INV_X1    g209(.A(G148gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n398_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n396_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n388_), .A2(KEYINPUT87), .A3(new_n398_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n415_), .A3(new_n395_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n392_), .B1(new_n416_), .B2(new_n393_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n391_), .B1(new_n408_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(KEYINPUT90), .B(new_n391_), .C1(new_n408_), .C2(new_n417_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n374_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n389_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n393_), .B1(new_n400_), .B2(new_n406_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT89), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n426_), .B2(new_n407_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n375_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n423_), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G85gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT0), .B(G57gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  AND2_X1   g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n420_), .A2(new_n435_), .A3(new_n374_), .A4(new_n421_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT102), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n422_), .A2(KEYINPUT4), .A3(new_n428_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n423_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n434_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n429_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n438_), .A2(new_n439_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n427_), .A2(KEYINPUT90), .ZN(new_n444_));
  AOI211_X1 g243(.A(new_n419_), .B(new_n424_), .C1(new_n426_), .C2(new_n407_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(KEYINPUT102), .A3(new_n435_), .A4(new_n374_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT102), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n436_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n442_), .B1(new_n443_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n441_), .B1(new_n451_), .B2(new_n433_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G22gat), .B(G50gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n454_), .B(KEYINPUT91), .Z(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n420_), .A2(new_n421_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  AOI211_X1 g259(.A(KEYINPUT29), .B(new_n456_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n455_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n456_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n455_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n458_), .A2(new_n459_), .A3(new_n457_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G78gat), .B(G106gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n462_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(KEYINPUT98), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G197gat), .A2(G204gat), .ZN(new_n474_));
  INV_X1    g273(.A(G197gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT93), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(G197gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n474_), .B1(new_n479_), .B2(G204gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT21), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G211gat), .B(G218gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT96), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G218gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n485_), .A2(G211gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(G211gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT96), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n480_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT97), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n480_), .A2(new_n484_), .A3(KEYINPUT97), .A4(new_n488_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n482_), .B1(new_n480_), .B2(KEYINPUT21), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n475_), .A2(G204gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(G204gat), .B1(new_n476_), .B2(new_n478_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AOI211_X1 g297(.A(KEYINPUT94), .B(G204gat), .C1(new_n476_), .C2(new_n478_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT21), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n494_), .B1(new_n500_), .B2(KEYINPUT95), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(KEYINPUT21), .C1(new_n498_), .C2(new_n499_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n493_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(G228gat), .A2(G233gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT99), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n427_), .A2(new_n459_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n505_), .B1(new_n509_), .B2(new_n504_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n507_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n470_), .A2(new_n473_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(new_n510_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT99), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n507_), .A2(new_n510_), .A3(new_n508_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n460_), .A2(new_n461_), .A3(new_n455_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n465_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n471_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n462_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n518_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n453_), .B1(new_n514_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G226gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n529_));
  NOR2_X1   g328(.A1(G183gat), .A2(G190gat), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n332_), .B1(new_n336_), .B2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n329_), .A2(new_n345_), .A3(new_n341_), .A4(new_n339_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n529_), .B1(new_n504_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT105), .ZN(new_n536_));
  INV_X1    g335(.A(new_n348_), .ZN(new_n537_));
  OAI22_X1  g336(.A1(new_n535_), .A2(new_n536_), .B1(new_n537_), .B2(new_n504_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n535_), .A2(new_n536_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n528_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n501_), .A2(new_n503_), .ZN(new_n541_));
  OAI211_X1 g340(.A(KEYINPUT101), .B(new_n533_), .C1(new_n541_), .C2(new_n493_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n529_), .B1(new_n504_), .B2(new_n537_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT101), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n504_), .B2(new_n534_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n540_), .B1(new_n528_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G8gat), .B(G36gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT18), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G64gat), .B(G92gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n528_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n504_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n528_), .B1(new_n555_), .B2(new_n348_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n535_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n554_), .A2(new_n551_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT27), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n552_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n551_), .A3(new_n557_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n559_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT106), .B1(new_n524_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n513_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n521_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n452_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n553_), .A2(new_n560_), .B1(new_n565_), .B2(new_n559_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT106), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n514_), .A2(new_n523_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n551_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n558_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n422_), .A2(new_n428_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n423_), .B1(new_n580_), .B2(KEYINPUT103), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT103), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n422_), .A2(new_n582_), .A3(new_n428_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n433_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n438_), .A2(new_n423_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n584_), .B(new_n585_), .C1(new_n437_), .C2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n429_), .A2(new_n433_), .ZN(new_n588_));
  AOI211_X1 g387(.A(KEYINPUT33), .B(new_n588_), .C1(new_n443_), .C2(new_n450_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n436_), .A2(new_n448_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n436_), .A2(new_n448_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n439_), .B(new_n438_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n593_), .B2(new_n434_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n579_), .B(new_n587_), .C1(new_n589_), .C2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT104), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n551_), .A2(KEYINPUT32), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n562_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n547_), .B2(new_n597_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n595_), .A2(new_n596_), .B1(new_n452_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n441_), .A2(KEYINPUT33), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n593_), .A2(new_n590_), .A3(new_n434_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n603_), .A2(KEYINPUT104), .A3(new_n579_), .A4(new_n587_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n577_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  OAI211_X1 g404(.A(KEYINPUT107), .B(new_n376_), .C1(new_n575_), .C2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n371_), .B(new_n374_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n576_), .A2(new_n572_), .A3(KEYINPUT108), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT108), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n577_), .B2(new_n567_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n607_), .A2(new_n608_), .A3(new_n610_), .A4(new_n453_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n589_), .A2(new_n594_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n585_), .B1(new_n437_), .B2(new_n586_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n581_), .A2(new_n583_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n563_), .B(new_n564_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n596_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n599_), .A2(new_n452_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n604_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n576_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n568_), .A3(new_n574_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT107), .B1(new_n621_), .B2(new_n376_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n612_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n286_), .B(KEYINPUT77), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n267_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(G229gat), .A3(G233gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT78), .Z(new_n627_));
  OR2_X1    g426(.A1(new_n624_), .A2(new_n267_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n267_), .A2(new_n289_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT79), .Z(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G113gat), .B(G141gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT80), .ZN(new_n635_));
  XOR2_X1   g434(.A(G169gat), .B(G197gat), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n633_), .B(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n623_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n321_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(new_n452_), .A3(new_n261_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n643_));
  OAI21_X1  g442(.A(new_n376_), .B1(new_n575_), .B2(new_n605_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n611_), .A3(new_n606_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n259_), .A2(new_n638_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n282_), .A2(new_n312_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n452_), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n642_), .A2(new_n643_), .B1(G1gat), .B2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n652_), .B1(new_n642_), .B2(new_n643_), .ZN(G1324gat));
  NAND3_X1  g452(.A1(new_n641_), .A2(new_n262_), .A3(new_n567_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n567_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G8gat), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(KEYINPUT39), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(KEYINPUT39), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g459(.A1(new_n650_), .A2(new_n607_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G15gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT41), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n640_), .A2(G15gat), .A3(new_n376_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n650_), .B2(new_n577_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT42), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n641_), .A2(new_n666_), .A3(new_n577_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n282_), .A2(new_n312_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n259_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n639_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT114), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT114), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n639_), .A2(new_n675_), .A3(new_n672_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n452_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n314_), .A2(new_n317_), .A3(KEYINPUT111), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT111), .B1(new_n314_), .B2(new_n317_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n612_), .B2(new_n622_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n319_), .A2(KEYINPUT43), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n682_), .A2(new_n684_), .B1(new_n647_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n648_), .A2(new_n282_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n693_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n683_), .B1(new_n647_), .B2(new_n681_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n319_), .A2(KEYINPUT43), .ZN(new_n696_));
  INV_X1    g495(.A(new_n612_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n646_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT112), .B(new_n689_), .C1(new_n695_), .C2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n694_), .A2(new_n691_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT113), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n694_), .A2(KEYINPUT113), .A3(new_n699_), .A4(new_n691_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n692_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n452_), .A2(G29gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n678_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(G36gat), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n674_), .A2(new_n707_), .A3(new_n567_), .A4(new_n676_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n567_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n711_), .B2(new_n707_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n709_), .B(KEYINPUT46), .C1(new_n711_), .C2(new_n707_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  INV_X1    g515(.A(G43gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n376_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n692_), .B(new_n719_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G43gat), .B1(new_n677_), .B2(new_n607_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT47), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n704_), .A2(new_n718_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(new_n721_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n723_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n722_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n677_), .B2(new_n577_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n577_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n704_), .B2(new_n729_), .ZN(G1331gat));
  INV_X1    g529(.A(new_n638_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n623_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n260_), .A3(new_n649_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G57gat), .B1(new_n733_), .B2(new_n453_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n732_), .A2(new_n259_), .A3(new_n283_), .A4(new_n319_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n453_), .A2(G57gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n733_), .B2(new_n572_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n572_), .A2(G64gat), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT115), .Z(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n735_), .B2(new_n741_), .ZN(G1333gat));
  OAI21_X1  g541(.A(G71gat), .B1(new_n733_), .B2(new_n376_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT49), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n376_), .A2(G71gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n735_), .B2(new_n745_), .ZN(G1334gat));
  OAI21_X1  g545(.A(G78gat), .B1(new_n733_), .B2(new_n576_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(KEYINPUT50), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(G78gat), .C1(new_n733_), .C2(new_n576_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n576_), .A2(G78gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT116), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n748_), .A2(new_n751_), .B1(new_n735_), .B2(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT117), .Z(G1335gat));
  INV_X1    g554(.A(new_n259_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n756_), .A2(new_n283_), .A3(new_n731_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n687_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n453_), .ZN(new_n759_));
  AND4_X1   g558(.A1(new_n260_), .A2(new_n732_), .A3(new_n282_), .A4(new_n312_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT118), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n453_), .A2(G85gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n758_), .B2(new_n572_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n572_), .A2(G92gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n758_), .B2(new_n376_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n376_), .A2(new_n213_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n761_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n760_), .B(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(G106gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n577_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G106gat), .B1(new_n758_), .B2(new_n576_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(KEYINPUT52), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n776_), .A2(KEYINPUT52), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n775_), .B(new_n781_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  INV_X1    g582(.A(new_n633_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n631_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n628_), .A2(new_n629_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n637_), .B1(new_n625_), .B2(new_n631_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n784_), .A2(new_n637_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n255_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n245_), .A2(new_n246_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n245_), .A2(new_n790_), .A3(new_n246_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n205_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(new_n796_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n731_), .A2(new_n254_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n797_), .B2(KEYINPUT119), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n789_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  OR3_X1    g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n312_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n795_), .A2(new_n796_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n254_), .B(new_n788_), .C1(new_n807_), .C2(new_n797_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n319_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n808_), .A2(KEYINPUT120), .A3(new_n809_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n788_), .A2(new_n254_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n814_), .B2(KEYINPUT58), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n810_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n805_), .B1(new_n804_), .B2(new_n312_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n806_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n282_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n756_), .A2(new_n638_), .A3(new_n283_), .A4(new_n319_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT54), .Z(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n607_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT59), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n823_), .A2(new_n452_), .A3(new_n824_), .A4(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n821_), .B1(new_n818_), .B2(new_n282_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n824_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n828_), .A2(new_n453_), .A3(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n638_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n830_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n638_), .A2(G113gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1340gat));
  INV_X1    g635(.A(new_n260_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G120gat), .B1(new_n832_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT60), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n259_), .A2(new_n839_), .ZN(new_n840_));
  MUX2_X1   g639(.A(new_n840_), .B(new_n839_), .S(G120gat), .Z(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n834_), .B2(new_n841_), .ZN(G1341gat));
  OAI21_X1  g641(.A(G127gat), .B1(new_n832_), .B2(new_n282_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n282_), .A2(G127gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n834_), .B2(new_n844_), .ZN(G1342gat));
  OAI21_X1  g644(.A(G134gat), .B1(new_n832_), .B2(new_n319_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n316_), .A2(G134gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n834_), .B2(new_n847_), .ZN(G1343gat));
  NOR2_X1   g647(.A1(new_n828_), .A2(new_n453_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n607_), .A2(new_n576_), .A3(new_n567_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n731_), .A3(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n260_), .A3(new_n850_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g653(.A1(new_n849_), .A2(new_n283_), .A3(new_n850_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  AND2_X1   g656(.A1(new_n849_), .A2(new_n850_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G162gat), .B1(new_n858_), .B2(new_n312_), .ZN(new_n859_));
  INV_X1    g658(.A(G162gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n679_), .A2(new_n680_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n858_), .B2(new_n861_), .ZN(G1347gat));
  NOR2_X1   g661(.A1(new_n376_), .A2(new_n452_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n567_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n823_), .A2(new_n576_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n868_));
  AND2_X1   g667(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n867_), .B(new_n731_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n823_), .A2(new_n576_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n865_), .A2(new_n731_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT122), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G169gat), .B1(new_n871_), .B2(new_n874_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n875_), .A2(KEYINPUT62), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(KEYINPUT62), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n870_), .B1(new_n876_), .B2(new_n877_), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n867_), .B2(new_n259_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n864_), .B1(new_n871_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n823_), .A2(KEYINPUT123), .A3(new_n576_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n260_), .A2(G176gat), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .A4(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n880_), .B1(new_n828_), .B2(new_n577_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n886_), .A2(new_n883_), .A3(new_n865_), .A4(new_n884_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT124), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n879_), .B1(new_n885_), .B2(new_n888_), .ZN(G1349gat));
  NOR3_X1   g688(.A1(new_n866_), .A2(new_n337_), .A3(new_n282_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n881_), .A2(new_n283_), .A3(new_n883_), .ZN(new_n891_));
  INV_X1    g690(.A(G183gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n866_), .B2(new_n319_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n312_), .A2(new_n338_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n866_), .B2(new_n895_), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n607_), .A2(new_n572_), .A3(new_n524_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n823_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n638_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n475_), .ZN(G1352gat));
  AND2_X1   g699(.A1(new_n823_), .A2(new_n897_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n260_), .A3(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT126), .Z(new_n905_));
  XNOR2_X1  g704(.A(new_n903_), .B(new_n905_), .ZN(G1353gat));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AND2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n898_), .A2(new_n282_), .A3(new_n907_), .A4(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n901_), .A2(new_n283_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n907_), .ZN(G1354gat));
  NAND3_X1  g710(.A1(new_n901_), .A2(new_n485_), .A3(new_n312_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G218gat), .B1(new_n898_), .B2(new_n319_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT127), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n916_), .A3(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1355gat));
endmodule


