//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(KEYINPUT92), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G197gat), .B(G204gat), .Z(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(KEYINPUT91), .A3(KEYINPUT21), .ZN(new_n205_));
  XOR2_X1   g004(.A(G211gat), .B(G218gat), .Z(new_n206_));
  OAI22_X1  g005(.A1(new_n205_), .A2(new_n206_), .B1(KEYINPUT21), .B2(new_n204_), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(KEYINPUT1), .B2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(KEYINPUT1), .ZN(new_n216_));
  AOI211_X1 g015(.A(new_n211_), .B(new_n212_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT2), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT87), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n210_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT88), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT88), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n225_), .B(new_n210_), .C1(new_n220_), .C2(new_n222_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n212_), .A2(KEYINPUT3), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(G141gat), .B2(G148gat), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n227_), .A2(new_n229_), .B1(new_n211_), .B2(KEYINPUT2), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n224_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n214_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(new_n213_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n231_), .A2(KEYINPUT89), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT89), .B1(new_n231_), .B2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n218_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n209_), .B1(new_n236_), .B2(KEYINPUT29), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT28), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n231_), .A2(new_n233_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT89), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n231_), .A2(KEYINPUT89), .A3(new_n233_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n217_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n239_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n237_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G22gat), .B(G50gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n207_), .A2(new_n208_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n249_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT28), .B1(new_n236_), .B2(KEYINPUT29), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n244_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n247_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n248_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n255_));
  INV_X1    g054(.A(G228gat), .ZN(new_n256_));
  INV_X1    g055(.A(G233gat), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT90), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(KEYINPUT90), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n256_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G78gat), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n254_), .A2(new_n255_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n248_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n253_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n247_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n263_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n203_), .B1(new_n262_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n261_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n263_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n202_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G8gat), .B(G36gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT23), .ZN(new_n281_));
  INV_X1    g080(.A(G169gat), .ZN(new_n282_));
  INV_X1    g081(.A(G176gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n281_), .B1(KEYINPUT24), .B2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G169gat), .B(G176gat), .Z(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(KEYINPUT24), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288_));
  INV_X1    g087(.A(G183gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT84), .B(G183gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(new_n288_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G190gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(KEYINPUT85), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT85), .B1(new_n292_), .B2(new_n293_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n287_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n291_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n281_), .B1(new_n298_), .B2(G190gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G169gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n209_), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n281_), .B1(new_n284_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n286_), .A2(new_n304_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT25), .B(G183gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n293_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT94), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n311_), .A3(new_n308_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n305_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n281_), .B1(G183gat), .B2(G190gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n314_), .A2(new_n301_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n249_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n303_), .A2(new_n316_), .A3(KEYINPUT20), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT19), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(KEYINPUT95), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n297_), .A2(new_n302_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n249_), .ZN(new_n322_));
  OR3_X1    g121(.A1(new_n313_), .A2(new_n249_), .A3(new_n315_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n319_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(KEYINPUT20), .A4(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT95), .B1(new_n317_), .B2(new_n319_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n279_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n317_), .A2(new_n319_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT95), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n279_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n325_), .A4(new_n320_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n322_), .A2(new_n323_), .A3(KEYINPUT20), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n319_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n317_), .A2(new_n319_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n333_), .B(KEYINPUT27), .C1(new_n340_), .C2(new_n332_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n274_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G71gat), .B(G99gat), .ZN(new_n344_));
  INV_X1    g143(.A(G43gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n321_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n346_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n297_), .A2(new_n302_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(G15gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT30), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT31), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n347_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n355_));
  OR3_X1    g154(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT86), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G113gat), .B(G120gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT86), .B1(new_n354_), .B2(new_n355_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n356_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G85gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n236_), .A2(new_n370_), .A3(new_n359_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT97), .ZN(new_n375_));
  INV_X1    g174(.A(new_n359_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT98), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n375_), .B(new_n376_), .C1(new_n236_), .C2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT97), .B1(new_n244_), .B2(KEYINPUT98), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n359_), .B1(new_n236_), .B2(new_n375_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n374_), .B1(new_n381_), .B2(KEYINPUT4), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n376_), .B1(new_n244_), .B2(KEYINPUT97), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n375_), .B1(new_n236_), .B2(new_n377_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n373_), .B1(new_n385_), .B2(new_n378_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n369_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n372_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n370_), .B1(new_n385_), .B2(new_n378_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n388_), .B(new_n368_), .C1(new_n389_), .C2(new_n374_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n364_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n343_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n336_), .A2(new_n390_), .A3(new_n387_), .A4(new_n341_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n363_), .B1(new_n274_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT99), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n382_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n369_), .B1(new_n381_), .B2(new_n372_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT99), .A3(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n372_), .B1(new_n381_), .B2(KEYINPUT101), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(KEYINPUT101), .B2(new_n381_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n381_), .A2(KEYINPUT4), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n371_), .A2(new_n372_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n368_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n334_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n398_), .A2(KEYINPUT33), .A3(new_n399_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n402_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n326_), .A2(new_n327_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n391_), .A2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n410_), .A2(new_n273_), .A3(new_n270_), .A4(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n395_), .A2(new_n416_), .A3(KEYINPUT102), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT102), .B1(new_n395_), .B2(new_n416_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n393_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G141gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G169gat), .B(G197gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  NOR2_X1   g221(.A1(new_n422_), .A2(KEYINPUT82), .ZN(new_n423_));
  XOR2_X1   g222(.A(G29gat), .B(G36gat), .Z(new_n424_));
  XOR2_X1   g223(.A(G43gat), .B(G50gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT15), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT74), .B(G1gat), .ZN(new_n428_));
  INV_X1    g227(.A(G8gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT14), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G15gat), .B(G22gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G1gat), .B(G8gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n435_));
  INV_X1    g234(.A(new_n433_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n430_), .A2(new_n436_), .A3(new_n431_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n435_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n437_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n436_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n427_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n443_), .B(KEYINPUT81), .Z(new_n444_));
  INV_X1    g243(.A(new_n426_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n442_), .B2(new_n438_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G229gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n442_), .A2(new_n445_), .A3(new_n438_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT79), .B1(new_n453_), .B2(new_n446_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n446_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n452_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n451_), .B1(new_n458_), .B2(new_n448_), .ZN(new_n459_));
  AOI211_X1 g258(.A(KEYINPUT80), .B(new_n447_), .C1(new_n454_), .C2(new_n457_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n450_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT83), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n450_), .B(new_n463_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n423_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n423_), .A3(new_n464_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n419_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G85gat), .B(G92gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  INV_X1    g271(.A(G106gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  AOI211_X1 g281(.A(KEYINPUT8), .B(new_n470_), .C1(new_n477_), .C2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n481_), .A3(KEYINPUT66), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n477_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n470_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT8), .B1(new_n490_), .B2(KEYINPUT67), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT66), .B1(new_n479_), .B2(new_n481_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(new_n476_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n470_), .B1(new_n493_), .B2(new_n487_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT67), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n484_), .B1(new_n491_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n470_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n499_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n482_), .ZN(new_n502_));
  XOR2_X1   g301(.A(KEYINPUT10), .B(G99gat), .Z(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n473_), .B2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n427_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT34), .ZN(new_n509_));
  OAI221_X1 g308(.A(new_n507_), .B1(KEYINPUT35), .B2(new_n509_), .C1(new_n445_), .C2(new_n506_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(KEYINPUT35), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G190gat), .B(G218gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G134gat), .B(G162gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(KEYINPUT36), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n515_), .B(KEYINPUT36), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT73), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT37), .ZN(new_n521_));
  INV_X1    g320(.A(new_n512_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n518_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n517_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT13), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G57gat), .B(G64gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G71gat), .B(G78gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT11), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n528_), .A2(KEYINPUT11), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(new_n529_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n528_), .A2(KEYINPUT11), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n530_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n506_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n490_), .A2(KEYINPUT67), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n483_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n505_), .ZN(new_n541_));
  OAI211_X1 g340(.A(KEYINPUT12), .B(new_n535_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT68), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n506_), .A2(new_n544_), .A3(KEYINPUT12), .A4(new_n535_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n536_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n534_), .B1(new_n497_), .B2(new_n505_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n548_), .B2(KEYINPUT12), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n538_), .A2(new_n539_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n541_), .B1(new_n551_), .B2(new_n484_), .ZN(new_n552_));
  OAI211_X1 g351(.A(KEYINPUT69), .B(new_n550_), .C1(new_n552_), .C2(new_n534_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT64), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n546_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n536_), .B2(new_n548_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G120gat), .B(G148gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT71), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT72), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n561_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n558_), .A2(new_n559_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n527_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(KEYINPUT13), .A3(new_n568_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n442_), .A2(new_n438_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT77), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(new_n535_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n535_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G127gat), .B(G155gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT16), .ZN(new_n584_));
  XOR2_X1   g383(.A(G183gat), .B(G211gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT78), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n586_), .B(KEYINPUT17), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n580_), .A2(new_n581_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n526_), .A2(new_n575_), .A3(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n469_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n391_), .A3(new_n428_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT103), .Z(new_n600_));
  INV_X1    g399(.A(new_n393_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n402_), .A2(new_n409_), .A3(new_n408_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n270_), .A2(new_n415_), .A3(new_n273_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n271_), .A2(new_n272_), .A3(new_n202_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n202_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n394_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n364_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n602_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n395_), .A2(new_n416_), .A3(KEYINPUT102), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n601_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n523_), .A2(new_n517_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n575_), .A2(KEYINPUT104), .A3(new_n468_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n617_));
  INV_X1    g416(.A(new_n467_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n465_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n619_), .B2(new_n574_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n616_), .A2(new_n620_), .A3(new_n594_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n615_), .A2(new_n391_), .A3(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n597_), .A2(new_n598_), .B1(G1gat), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n600_), .A2(new_n623_), .ZN(G1324gat));
  INV_X1    g423(.A(KEYINPUT40), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT106), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n419_), .A2(new_n621_), .A3(new_n342_), .A4(new_n613_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT105), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G8gat), .B1(new_n627_), .B2(KEYINPUT105), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n627_), .A2(KEYINPUT105), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n632_), .A2(KEYINPUT106), .A3(G8gat), .A4(new_n628_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n631_), .A2(new_n633_), .A3(KEYINPUT39), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n626_), .B(new_n635_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n596_), .A2(new_n429_), .A3(new_n342_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n625_), .B1(new_n634_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n631_), .A2(new_n633_), .A3(KEYINPUT39), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n640_), .A2(KEYINPUT40), .A3(new_n636_), .A4(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(G1325gat));
  NAND3_X1  g441(.A1(new_n615_), .A2(new_n363_), .A3(new_n621_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT41), .B1(new_n643_), .B2(G15gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n596_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n364_), .A2(G15gat), .ZN(new_n647_));
  OAI22_X1  g446(.A1(new_n644_), .A2(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT107), .ZN(G1326gat));
  NAND3_X1  g448(.A1(new_n615_), .A2(new_n274_), .A3(new_n621_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G22gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  INV_X1    g451(.A(new_n274_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(G22gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(new_n646_), .B2(new_n654_), .ZN(G1327gat));
  INV_X1    g454(.A(new_n526_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n419_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n594_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n616_), .A2(new_n620_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n419_), .A2(KEYINPUT43), .A3(new_n656_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n658_), .B1(new_n612_), .B2(new_n526_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(new_n663_), .A3(new_n593_), .A4(new_n660_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n661_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n664_), .A2(new_n667_), .A3(G29gat), .A4(new_n391_), .ZN(new_n668_));
  INV_X1    g467(.A(G29gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n612_), .A2(new_n619_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n594_), .A2(new_n613_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n574_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n391_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n669_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n668_), .A2(new_n676_), .ZN(G1328gat));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n664_), .A2(new_n667_), .A3(new_n342_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  INV_X1    g483(.A(new_n342_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n670_), .A2(new_n684_), .A3(new_n673_), .A4(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n419_), .A2(new_n468_), .A3(new_n673_), .A4(new_n686_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT45), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n678_), .A2(new_n679_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n681_), .B1(new_n683_), .B2(new_n693_), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n680_), .B(new_n692_), .C1(new_n682_), .C2(G36gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1329gat));
  NAND4_X1  g495(.A1(new_n664_), .A2(new_n667_), .A3(G43gat), .A4(new_n363_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n345_), .B1(new_n674_), .B2(new_n364_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g499(.A1(new_n664_), .A2(new_n667_), .A3(G50gat), .A4(new_n274_), .ZN(new_n701_));
  INV_X1    g500(.A(G50gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n674_), .B2(new_n653_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1331gat));
  NOR3_X1   g503(.A1(new_n575_), .A2(new_n468_), .A3(new_n593_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n615_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(G57gat), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n675_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT112), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n526_), .A2(new_n594_), .A3(new_n574_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT110), .Z(new_n711_));
  NOR2_X1   g510(.A1(new_n612_), .A2(new_n468_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n391_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n713_), .A2(KEYINPUT111), .A3(new_n707_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT111), .B1(new_n713_), .B2(new_n707_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n709_), .A2(new_n714_), .A3(new_n715_), .ZN(G1332gat));
  OAI21_X1  g515(.A(G64gat), .B1(new_n706_), .B2(new_n685_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT48), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n711_), .A2(new_n712_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n685_), .A2(G64gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(G1333gat));
  OR3_X1    g520(.A1(new_n719_), .A2(G71gat), .A3(new_n364_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n615_), .A2(new_n363_), .A3(new_n705_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G71gat), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT49), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(KEYINPUT49), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1334gat));
  OAI21_X1  g528(.A(G78gat), .B1(new_n706_), .B2(new_n653_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT50), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n653_), .A2(G78gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n719_), .B2(new_n732_), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n575_), .A2(new_n468_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n665_), .A2(new_n663_), .A3(new_n593_), .A4(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n736_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n391_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G85gat), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n672_), .A2(new_n575_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n712_), .A2(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n675_), .A2(G85gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(G1336gat));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n342_), .A3(new_n738_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G92gat), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n685_), .A2(G92gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n742_), .B2(new_n747_), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n735_), .B2(new_n364_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n363_), .A2(new_n503_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n742_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g551(.A1(new_n712_), .A2(new_n473_), .A3(new_n274_), .A4(new_n741_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n659_), .A2(new_n274_), .A3(new_n663_), .A4(new_n734_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G106gat), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n754_), .B(G106gat), .C1(new_n735_), .C2(new_n653_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n753_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n753_), .C1(new_n756_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764_));
  INV_X1    g563(.A(new_n595_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n619_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n595_), .A2(KEYINPUT54), .A3(new_n468_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n468_), .A2(new_n568_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n557_), .B1(new_n546_), .B2(new_n554_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n558_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n546_), .A2(new_n554_), .A3(KEYINPUT55), .A4(new_n557_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n566_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n567_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT115), .B1(new_n779_), .B2(KEYINPUT56), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n779_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT116), .B1(new_n779_), .B2(KEYINPUT56), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n769_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n448_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n786_));
  OR3_X1    g585(.A1(new_n786_), .A2(KEYINPUT117), .A3(new_n422_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n444_), .A2(new_n455_), .A3(new_n448_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT117), .B1(new_n786_), .B2(new_n422_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n450_), .B(new_n422_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n572_), .B2(new_n568_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT57), .B(new_n613_), .C1(new_n785_), .C2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n779_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n778_), .A2(new_n798_), .A3(new_n780_), .A4(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n619_), .A2(new_n569_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n793_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n795_), .B1(new_n802_), .B2(new_n614_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n792_), .B2(new_n569_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n790_), .A2(KEYINPUT118), .A3(new_n568_), .A4(new_n791_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n779_), .A2(KEYINPUT56), .ZN(new_n808_));
  INV_X1    g607(.A(new_n796_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n807_), .B(KEYINPUT58), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n656_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n794_), .A2(new_n803_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n768_), .B1(new_n815_), .B2(new_n593_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n343_), .A2(new_n391_), .A3(new_n363_), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT119), .Z(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(G113gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n468_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(KEYINPUT59), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n619_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n822_), .B1(new_n826_), .B2(new_n821_), .ZN(G1340gat));
  INV_X1    g626(.A(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n575_), .B2(KEYINPUT60), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n820_), .B(new_n829_), .C1(KEYINPUT60), .C2(new_n828_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n575_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n828_), .ZN(G1341gat));
  INV_X1    g631(.A(G127gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n820_), .A2(new_n833_), .A3(new_n594_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n593_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n833_), .ZN(G1342gat));
  NOR3_X1   g635(.A1(new_n816_), .A2(new_n613_), .A3(new_n819_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(KEYINPUT120), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n837_), .B2(G134gat), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n823_), .A2(new_n825_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n526_), .A2(new_n839_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT121), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n840_), .A2(new_n842_), .B1(new_n843_), .B2(new_n845_), .ZN(G1343gat));
  NAND2_X1  g645(.A1(new_n815_), .A2(new_n593_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n768_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NOR4_X1   g648(.A1(new_n653_), .A2(new_n675_), .A3(new_n342_), .A4(new_n363_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n468_), .A3(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n850_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n575_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT122), .B(G148gat), .Z(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1345gat));
  NAND3_X1  g655(.A1(new_n849_), .A2(new_n594_), .A3(new_n850_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  INV_X1    g658(.A(G162gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n853_), .A2(new_n860_), .A3(new_n526_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n849_), .A2(new_n614_), .A3(new_n850_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT123), .B1(new_n862_), .B2(G162gat), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n864_), .B(new_n860_), .C1(new_n853_), .C2(new_n613_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n861_), .B1(new_n863_), .B2(new_n865_), .ZN(G1347gat));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n653_), .A2(new_n342_), .A3(new_n392_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n849_), .A2(new_n867_), .A3(new_n468_), .A4(new_n869_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n816_), .A2(KEYINPUT22), .A3(new_n619_), .A4(new_n868_), .ZN(new_n871_));
  OAI211_X1 g670(.A(G169gat), .B(new_n870_), .C1(new_n871_), .C2(new_n867_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n816_), .A2(new_n868_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT22), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n468_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT62), .A3(new_n282_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n872_), .A2(new_n876_), .ZN(G1348gat));
  NOR3_X1   g676(.A1(new_n816_), .A2(new_n575_), .A3(new_n868_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n283_), .A2(KEYINPUT124), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n283_), .A2(KEYINPUT124), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n878_), .B2(new_n880_), .ZN(G1349gat));
  NOR3_X1   g681(.A1(new_n816_), .A2(new_n593_), .A3(new_n868_), .ZN(new_n883_));
  MUX2_X1   g682(.A(new_n298_), .B(new_n307_), .S(new_n883_), .Z(G1350gat));
  NAND2_X1  g683(.A1(new_n614_), .A2(new_n293_), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT125), .Z(new_n886_));
  NAND2_X1  g685(.A1(new_n873_), .A2(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n816_), .A2(new_n526_), .A3(new_n868_), .ZN(new_n888_));
  INV_X1    g687(.A(G190gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1351gat));
  NAND3_X1  g689(.A1(new_n364_), .A2(new_n675_), .A3(new_n342_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n816_), .A2(new_n653_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n468_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g693(.A(new_n575_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n892_), .A2(new_n895_), .ZN(new_n896_));
  OR2_X1    g695(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1353gat));
  NAND2_X1  g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n594_), .A3(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT127), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n903_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n892_), .A2(new_n594_), .A3(new_n902_), .A4(new_n899_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1354gat));
  INV_X1    g705(.A(G218gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n892_), .A2(new_n907_), .A3(new_n614_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n892_), .A2(new_n656_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1355gat));
endmodule


