//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n958_, new_n959_,
    new_n960_, new_n962_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n991_, new_n992_, new_n993_;
  INV_X1    g000(.A(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT6), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G85gat), .B(G92gat), .Z(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(KEYINPUT9), .B2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT10), .B(G99gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(new_n203_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n210_), .B(new_n212_), .C1(KEYINPUT9), .C2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(new_n202_), .A3(new_n203_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n215_), .B(new_n209_), .C1(new_n208_), .C2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n218_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT64), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n217_), .A2(new_n224_), .A3(new_n218_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n207_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n215_), .B1(new_n226_), .B2(new_n209_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n220_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n209_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n219_), .A2(KEYINPUT64), .B1(new_n204_), .B2(new_n206_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(new_n225_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n232_), .A2(KEYINPUT65), .A3(new_n215_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n214_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G29gat), .B(G36gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G43gat), .B(G50gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT15), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(new_n232_), .B2(new_n215_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n227_), .A2(new_n228_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n220_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(new_n214_), .A3(new_n237_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G232gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT34), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT35), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n240_), .A2(new_n244_), .A3(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n247_), .A2(new_n248_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n240_), .A2(new_n253_), .A3(new_n244_), .A4(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G190gat), .B(G218gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G134gat), .B(G162gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT36), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT67), .B(KEYINPUT36), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n252_), .A2(new_n254_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(KEYINPUT37), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n259_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n255_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n267_), .B2(new_n255_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n263_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT37), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n265_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G15gat), .B(G22gat), .ZN(new_n273_));
  INV_X1    g072(.A(G1gat), .ZN(new_n274_));
  INV_X1    g073(.A(G8gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT14), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G1gat), .B(G8gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT70), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT70), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT71), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n285_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G57gat), .B(G64gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT66), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G71gat), .B(G78gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n290_), .B(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n292_), .A2(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n288_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n288_), .A2(new_n299_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G155gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT17), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n302_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n302_), .A2(new_n309_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(KEYINPUT73), .B2(new_n311_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n272_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT74), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT86), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G155gat), .A3(G162gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n325_), .B2(KEYINPUT1), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(new_n324_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT87), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT87), .A4(new_n327_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n326_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT85), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G141gat), .A3(G148gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G141gat), .ZN(new_n338_));
  INV_X1    g137(.A(G148gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n332_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n334_), .A2(new_n336_), .A3(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n338_), .A2(new_n339_), .A3(KEYINPUT3), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(G141gat), .B2(G148gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n320_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT88), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n350_), .A2(KEYINPUT88), .A3(new_n351_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n341_), .B(new_n342_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT89), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n351_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT88), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n350_), .A2(KEYINPUT88), .A3(new_n351_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(KEYINPUT89), .A3(new_n342_), .A4(new_n341_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G22gat), .B(G50gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT28), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n356_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(G228gat), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n341_), .B1(new_n353_), .B2(new_n352_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(KEYINPUT92), .A2(G197gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(KEYINPUT92), .A2(G197gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n375_), .B1(new_n378_), .B2(G204gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G211gat), .B(G218gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT21), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G204gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n376_), .A2(new_n384_), .A3(new_n377_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n381_), .B1(G197gat), .B2(G204gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n380_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n377_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(KEYINPUT92), .A2(G197gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(G204gat), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n375_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT21), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n383_), .B1(new_n388_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT91), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n372_), .B1(new_n374_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n372_), .ZN(new_n398_));
  AOI211_X1 g197(.A(new_n398_), .B(new_n395_), .C1(new_n373_), .C2(KEYINPUT29), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n368_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n342_), .B1(new_n361_), .B2(new_n341_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n401_), .B2(new_n395_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n374_), .A2(new_n372_), .A3(new_n396_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n368_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n367_), .A2(new_n400_), .A3(KEYINPUT93), .A4(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT93), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n409_), .A2(new_n367_), .B1(new_n400_), .B2(new_n405_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G127gat), .B(G134gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G113gat), .B(G120gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT84), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT31), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n414_), .A2(KEYINPUT84), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(KEYINPUT84), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT31), .A3(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(G15gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT30), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n426_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n417_), .A2(new_n418_), .A3(new_n421_), .A4(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT79), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT77), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n433_), .A2(KEYINPUT78), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT25), .B(G183gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT26), .B(G190gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n437_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT78), .B1(new_n445_), .B2(new_n433_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n431_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n436_), .A2(new_n437_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n432_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n450_), .A2(KEYINPUT79), .A3(new_n438_), .A4(new_n441_), .ZN(new_n451_));
  AND3_X1   g250(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT24), .ZN(new_n455_));
  INV_X1    g254(.A(G169gat), .ZN(new_n456_));
  INV_X1    g255(.A(G176gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT80), .B1(new_n454_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G183gat), .A2(G190gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT23), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n463_));
  AND4_X1   g262(.A1(KEYINPUT80), .A2(new_n458_), .A3(new_n462_), .A4(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n447_), .A2(new_n451_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n456_), .B2(KEYINPUT22), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT22), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT81), .A3(G169gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n456_), .A2(KEYINPUT22), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n468_), .A2(new_n470_), .A3(new_n457_), .A4(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n472_), .A2(KEYINPUT82), .A3(new_n445_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT82), .B1(new_n472_), .B2(new_n445_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G183gat), .A2(G190gat), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n452_), .A2(new_n453_), .A3(new_n475_), .ZN(new_n476_));
  OR3_X1    g275(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n466_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G71gat), .B(G99gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G43gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n478_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n430_), .B(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n411_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G226gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT19), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n440_), .B(KEYINPUT94), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n439_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n454_), .A2(new_n458_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n434_), .B2(new_n433_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n476_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT22), .B(G169gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n457_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n495_), .A3(new_n445_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT20), .B1(new_n497_), .B2(new_n394_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT95), .B1(new_n478_), .B2(new_n394_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT95), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n387_), .A2(new_n380_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n391_), .A2(new_n392_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n381_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n502_), .A2(new_n504_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n501_), .B(new_n505_), .C1(new_n466_), .C2(new_n477_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n487_), .B(new_n499_), .C1(new_n500_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n497_), .B2(new_n394_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(new_n394_), .B2(new_n478_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n486_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G8gat), .B(G36gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT18), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G64gat), .B(G92gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  AND3_X1   g314(.A1(new_n507_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT96), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n507_), .A2(new_n511_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n515_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT96), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n507_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G29gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(G85gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT0), .B(G57gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G225gat), .A2(G233gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n341_), .B(KEYINPUT97), .C1(new_n352_), .C2(new_n353_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n414_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n414_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n361_), .A2(KEYINPUT97), .A3(new_n341_), .A4(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n532_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n359_), .A2(new_n360_), .B1(new_n332_), .B2(new_n340_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n538_), .A2(KEYINPUT4), .A3(new_n414_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n531_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n534_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n529_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n542_), .A2(new_n543_), .A3(KEYINPUT33), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n542_), .B2(KEYINPUT33), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n518_), .B(new_n524_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n535_), .B1(new_n538_), .B2(KEYINPUT97), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n533_), .A2(new_n414_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT4), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n539_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n530_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n534_), .A2(new_n536_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n528_), .B1(new_n552_), .B2(new_n531_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT100), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT100), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n530_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n541_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n528_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT99), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT99), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n542_), .A2(new_n564_), .A3(KEYINPUT33), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n558_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n546_), .A2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n509_), .B(new_n487_), .C1(new_n394_), .C2(new_n478_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n451_), .A2(new_n465_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(new_n447_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n501_), .B1(new_n571_), .B2(new_n505_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n478_), .A2(KEYINPUT95), .A3(new_n394_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n498_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n568_), .B1(new_n574_), .B2(new_n487_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n515_), .A2(KEYINPUT32), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n507_), .A2(new_n511_), .A3(new_n576_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n540_), .A2(new_n541_), .A3(new_n529_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n578_), .B(new_n579_), .C1(new_n581_), .C2(new_n542_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n561_), .A2(new_n580_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n585_), .A2(KEYINPUT101), .A3(new_n579_), .A4(new_n578_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n484_), .B1(new_n567_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n483_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n409_), .A2(new_n367_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n400_), .A2(new_n405_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n481_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n481_), .B1(new_n429_), .B2(new_n427_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(new_n595_), .A3(new_n406_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n589_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT27), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n521_), .A2(new_n523_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n523_), .A2(KEYINPUT27), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n515_), .B(KEYINPUT102), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n575_), .A2(new_n601_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n598_), .A2(new_n599_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n585_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n597_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n588_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT5), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(KEYINPUT12), .ZN(new_n612_));
  INV_X1    g411(.A(new_n299_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n234_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n243_), .A2(new_n214_), .A3(new_n299_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n299_), .B1(new_n243_), .B2(new_n214_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(KEYINPUT12), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n616_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n611_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n615_), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT12), .B1(new_n624_), .B2(new_n617_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n614_), .A2(new_n612_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n619_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n622_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n611_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT13), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n623_), .A2(KEYINPUT13), .A3(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT75), .ZN(new_n637_));
  INV_X1    g436(.A(new_n284_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n237_), .B1(new_n638_), .B2(new_n282_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n237_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n283_), .A2(new_n640_), .A3(new_n284_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n638_), .A2(new_n237_), .A3(new_n282_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(KEYINPUT75), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n636_), .B1(new_n642_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT76), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n643_), .B1(new_n238_), .B2(new_n285_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n636_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT76), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n646_), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G113gat), .B(G141gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G169gat), .B(G197gat), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n653_), .B(new_n654_), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n652_), .B(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n635_), .A2(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n319_), .A2(new_n607_), .A3(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n274_), .A3(new_n585_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT38), .Z(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n317_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n607_), .A2(new_n663_), .A3(new_n270_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n584_), .B(new_n586_), .C1(new_n546_), .C2(new_n566_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n605_), .B1(new_n665_), .B2(new_n484_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n270_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT103), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n662_), .B1(new_n664_), .B2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n274_), .B1(new_n669_), .B2(new_n585_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n661_), .A2(new_n670_), .ZN(G1324gat));
  INV_X1    g470(.A(new_n603_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n659_), .A2(new_n275_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n669_), .A2(new_n672_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(G8gat), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT39), .B(new_n275_), .C1(new_n669_), .C2(new_n672_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1325gat));
  NAND3_X1  g479(.A1(new_n659_), .A2(new_n424_), .A3(new_n483_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n669_), .A2(new_n483_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT41), .B1(new_n682_), .B2(G15gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(new_n411_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(G22gat), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT104), .Z(new_n688_));
  NAND2_X1  g487(.A1(new_n659_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n669_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G22gat), .B1(new_n690_), .B2(new_n686_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(KEYINPUT42), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(KEYINPUT42), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(G1327gat));
  NOR2_X1   g493(.A1(new_n317_), .A2(new_n270_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n484_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n584_), .A2(new_n586_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n518_), .A2(new_n524_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT98), .B1(new_n561_), .B2(new_n562_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n542_), .A2(new_n543_), .A3(KEYINPUT33), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n561_), .A2(KEYINPUT99), .A3(new_n562_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n564_), .B1(new_n542_), .B2(KEYINPUT33), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n698_), .A2(new_n701_), .A3(new_n704_), .A4(new_n558_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n696_), .B1(new_n697_), .B2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n658_), .B(new_n695_), .C1(new_n706_), .C2(new_n605_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT106), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n607_), .A2(new_n709_), .A3(new_n658_), .A4(new_n695_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n604_), .A2(G29gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n666_), .B2(new_n272_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  INV_X1    g513(.A(new_n272_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n714_), .B(new_n715_), .C1(new_n706_), .C2(new_n605_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n658_), .A2(new_n316_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n721_), .B(new_n718_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n585_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n724_), .A2(KEYINPUT105), .A3(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT105), .B1(new_n724_), .B2(G29gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n712_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n603_), .A2(G36gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n708_), .A2(new_n710_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n708_), .A2(new_n710_), .A3(KEYINPUT45), .A4(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n714_), .B1(new_n607_), .B2(new_n715_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n666_), .A2(KEYINPUT43), .A3(new_n272_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n719_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n721_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n717_), .A2(KEYINPUT44), .A3(new_n719_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n672_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n734_), .B1(new_n740_), .B2(G36gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n728_), .B1(new_n741_), .B2(KEYINPUT107), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n743_));
  INV_X1    g542(.A(G36gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n723_), .B2(new_n672_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n743_), .B(KEYINPUT46), .C1(new_n745_), .C2(new_n734_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1329gat));
  NAND3_X1  g546(.A1(new_n723_), .A2(G43gat), .A3(new_n483_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n708_), .A2(new_n483_), .A3(new_n710_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT108), .B(G43gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(G1330gat));
  INV_X1    g553(.A(G50gat), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n686_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n708_), .A2(new_n411_), .A3(new_n710_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n723_), .A2(new_n756_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT110), .Z(G1331gat));
  AND2_X1   g558(.A1(new_n633_), .A2(new_n634_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n666_), .A2(new_n656_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n319_), .A2(new_n761_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n762_), .A2(G57gat), .A3(new_n604_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n760_), .A2(new_n656_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n317_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n664_), .B2(new_n668_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n585_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n763_), .B1(new_n767_), .B2(G57gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT111), .ZN(G1332gat));
  INV_X1    g568(.A(G64gat), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n319_), .A2(new_n761_), .A3(new_n770_), .A4(new_n672_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(new_n672_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(G64gat), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(G64gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(G1333gat));
  OR3_X1    g577(.A1(new_n762_), .A2(G71gat), .A3(new_n595_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n766_), .A2(new_n483_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G71gat), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT49), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(KEYINPUT49), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(G1334gat));
  OR3_X1    g583(.A1(new_n762_), .A2(G78gat), .A3(new_n686_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n766_), .A2(new_n411_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(G78gat), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G78gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(G1335gat));
  NAND3_X1  g589(.A1(new_n717_), .A2(new_n316_), .A3(new_n764_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791_), .B2(new_n604_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n761_), .A2(new_n695_), .ZN(new_n793_));
  OR3_X1    g592(.A1(new_n793_), .A2(G85gat), .A3(new_n604_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1336gat));
  INV_X1    g594(.A(G92gat), .ZN(new_n796_));
  OR3_X1    g595(.A1(new_n791_), .A2(new_n796_), .A3(new_n603_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n793_), .B2(new_n603_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n799_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n797_), .A2(new_n800_), .A3(new_n801_), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n791_), .B2(new_n595_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n483_), .A2(new_n211_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n793_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g605(.A1(new_n717_), .A2(new_n411_), .A3(new_n316_), .A4(new_n764_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n807_), .A2(new_n808_), .A3(G106gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n807_), .B2(G106gat), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n411_), .A2(new_n203_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n809_), .A2(new_n810_), .B1(new_n793_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g612(.A(new_n589_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n672_), .A2(new_n604_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n656_), .A2(new_n630_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n619_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n627_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n616_), .A2(new_n618_), .A3(new_n819_), .A4(new_n620_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n611_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n825_), .B(new_n629_), .C1(new_n820_), .C2(new_n822_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n817_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n650_), .B1(new_n642_), .B2(new_n645_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT116), .B1(new_n828_), .B2(new_n655_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n636_), .B1(new_n649_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n830_), .B2(new_n649_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n829_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n642_), .A2(new_n645_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n636_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836_));
  INV_X1    g635(.A(new_n655_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n833_), .A2(new_n838_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n631_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n631_), .B2(new_n839_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n827_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT57), .B1(new_n844_), .B2(new_n270_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n846_), .B(new_n667_), .C1(new_n827_), .C2(new_n843_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n839_), .A2(new_n630_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n272_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n620_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n621_), .B1(KEYINPUT55), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n611_), .B1(new_n854_), .B2(new_n821_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n825_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n611_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(KEYINPUT58), .A4(new_n849_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT58), .B(new_n849_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT119), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n852_), .A2(new_n860_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n317_), .B1(new_n848_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n265_), .B(new_n316_), .C1(new_n271_), .C2(new_n270_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n635_), .A2(new_n656_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AND4_X1   g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n317_), .A4(new_n272_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n814_), .B(new_n815_), .C1(new_n864_), .C2(new_n870_), .ZN(new_n871_));
  OR2_X1    g670(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n815_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n816_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n631_), .A2(new_n839_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT118), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n631_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n270_), .B1(new_n875_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n846_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n844_), .A2(KEYINPUT57), .A3(new_n270_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n863_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n316_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n870_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n874_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n814_), .A3(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n873_), .A2(new_n656_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G113gat), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n871_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n886_), .A2(KEYINPUT120), .A3(new_n814_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n657_), .A2(G113gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n890_), .A2(new_n895_), .ZN(G1340gat));
  NAND3_X1  g695(.A1(new_n873_), .A2(new_n635_), .A3(new_n888_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G120gat), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899_));
  AOI21_X1  g698(.A(G120gat), .B1(new_n635_), .B2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n899_), .B2(G120gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n892_), .A2(new_n893_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n902_), .ZN(G1341gat));
  AND2_X1   g702(.A1(new_n873_), .A2(new_n888_), .ZN(new_n904_));
  INV_X1    g703(.A(G127gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n316_), .A2(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT122), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n892_), .A2(new_n317_), .A3(new_n893_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n904_), .A2(new_n907_), .B1(new_n908_), .B2(new_n905_), .ZN(G1342gat));
  NAND3_X1  g708(.A1(new_n873_), .A2(new_n715_), .A3(new_n888_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G134gat), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n270_), .A2(G134gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n892_), .A2(new_n893_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1343gat));
  INV_X1    g713(.A(new_n596_), .ZN(new_n915_));
  AOI21_X1  g714(.A(KEYINPUT123), .B1(new_n886_), .B2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n870_), .B1(new_n883_), .B2(new_n316_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n917_), .A2(new_n918_), .A3(new_n596_), .A4(new_n874_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n656_), .B1(new_n916_), .B2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G141gat), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n338_), .B(new_n656_), .C1(new_n916_), .C2(new_n919_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1344gat));
  OAI21_X1  g722(.A(new_n635_), .B1(new_n916_), .B2(new_n919_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G148gat), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n339_), .B(new_n635_), .C1(new_n916_), .C2(new_n919_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1345gat));
  OAI21_X1  g726(.A(new_n317_), .B1(new_n916_), .B2(new_n919_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT61), .B(G155gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n929_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n317_), .B(new_n931_), .C1(new_n916_), .C2(new_n919_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1346gat));
  INV_X1    g732(.A(G162gat), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n934_), .B(new_n667_), .C1(new_n916_), .C2(new_n919_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n886_), .A2(new_n915_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n918_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n886_), .A2(KEYINPUT123), .A3(new_n915_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n272_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n935_), .B1(new_n939_), .B2(new_n934_), .ZN(G1347gat));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n884_), .A2(new_n885_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n603_), .A2(new_n585_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n483_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n686_), .A3(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n657_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n941_), .B1(new_n947_), .B2(new_n456_), .ZN(new_n948_));
  OAI211_X1 g747(.A(KEYINPUT62), .B(G169gat), .C1(new_n946_), .C2(new_n657_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n494_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n948_), .A2(new_n949_), .A3(new_n950_), .ZN(G1348gat));
  OR3_X1    g750(.A1(new_n917_), .A2(KEYINPUT124), .A3(new_n411_), .ZN(new_n952_));
  OAI21_X1  g751(.A(KEYINPUT124), .B1(new_n917_), .B2(new_n411_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n944_), .A2(new_n760_), .A3(new_n457_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n952_), .A2(new_n953_), .A3(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n457_), .B1(new_n946_), .B2(new_n760_), .ZN(new_n956_));
  AND2_X1   g755(.A1(new_n955_), .A2(new_n956_), .ZN(G1349gat));
  NOR3_X1   g756(.A1(new_n946_), .A2(new_n439_), .A3(new_n316_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n952_), .A2(new_n317_), .A3(new_n945_), .A4(new_n953_), .ZN(new_n959_));
  INV_X1    g758(.A(G183gat), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n958_), .B1(new_n959_), .B2(new_n960_), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n946_), .B2(new_n272_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n667_), .A2(new_n488_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(KEYINPUT125), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n962_), .B1(new_n946_), .B2(new_n964_), .ZN(G1351gat));
  NAND2_X1  g764(.A1(new_n943_), .A2(new_n915_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n942_), .A2(KEYINPUT126), .A3(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n969_), .B1(new_n917_), .B2(new_n966_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n970_), .ZN(new_n971_));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971_), .B2(new_n656_), .ZN(new_n972_));
  INV_X1    g771(.A(G197gat), .ZN(new_n973_));
  AOI211_X1 g772(.A(new_n973_), .B(new_n657_), .C1(new_n968_), .C2(new_n970_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n972_), .A2(new_n974_), .ZN(G1352gat));
  AOI21_X1  g774(.A(KEYINPUT126), .B1(new_n942_), .B2(new_n967_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n917_), .A2(new_n969_), .A3(new_n966_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n976_), .A2(new_n977_), .ZN(new_n978_));
  OAI21_X1  g777(.A(G204gat), .B1(new_n978_), .B2(new_n760_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n971_), .A2(new_n384_), .A3(new_n635_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1353gat));
  AOI21_X1  g780(.A(new_n316_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n982_), .B1(new_n976_), .B2(new_n977_), .ZN(new_n983_));
  OAI21_X1  g782(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n984_));
  NOR2_X1   g783(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n985_));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n985_), .A2(new_n986_), .ZN(new_n987_));
  NAND3_X1  g786(.A1(new_n983_), .A2(new_n984_), .A3(new_n987_), .ZN(new_n988_));
  NAND4_X1  g787(.A1(new_n971_), .A2(new_n986_), .A3(new_n982_), .A4(new_n985_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n988_), .A2(new_n989_), .ZN(G1354gat));
  OAI21_X1  g789(.A(G218gat), .B1(new_n978_), .B2(new_n272_), .ZN(new_n991_));
  INV_X1    g790(.A(G218gat), .ZN(new_n992_));
  NAND3_X1  g791(.A1(new_n971_), .A2(new_n992_), .A3(new_n667_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n991_), .A2(new_n993_), .ZN(G1355gat));
endmodule


