//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT3), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT2), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT91), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT91), .B1(new_n206_), .B2(new_n208_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n203_), .B(new_n204_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n202_), .B1(KEYINPUT1), .B2(new_n204_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(KEYINPUT1), .B2(new_n204_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n205_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n207_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G127gat), .B(G134gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G113gat), .B(G120gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n220_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT87), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n218_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n224_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(new_n221_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n213_), .A2(new_n217_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT4), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(new_n233_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G1gat), .B(G29gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G85gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G57gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n245_), .A3(new_n238_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT86), .Z(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G169gat), .ZN(new_n251_));
  INV_X1    g050(.A(G176gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT23), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT83), .B(G183gat), .Z(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(G190gat), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT85), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n250_), .A2(KEYINPUT24), .A3(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(new_n256_), .C1(KEYINPUT24), .C2(new_n261_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G190gat), .ZN(new_n264_));
  INV_X1    g063(.A(G183gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT25), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT84), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n264_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n257_), .B1(KEYINPUT84), .B2(new_n265_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(KEYINPUT25), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n259_), .B1(new_n263_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G43gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n271_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277_));
  INV_X1    g076(.A(G15gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT30), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n226_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n276_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n248_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G78gat), .B(G106gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT94), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT21), .ZN(new_n287_));
  XOR2_X1   g086(.A(G211gat), .B(G218gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(G197gat), .B(G204gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(KEYINPUT92), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(new_n288_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n288_), .B1(KEYINPUT92), .B2(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n287_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G228gat), .A2(G233gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n286_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(KEYINPUT94), .A3(new_n298_), .A4(new_n297_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n298_), .B1(new_n303_), .B2(new_n295_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n285_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI211_X1 g108(.A(new_n284_), .B(new_n306_), .C1(new_n302_), .C2(new_n304_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n213_), .A2(new_n300_), .A3(new_n217_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G22gat), .B(G50gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT28), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n312_), .B(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n309_), .A2(new_n311_), .A3(KEYINPUT95), .A4(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n306_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT95), .B1(new_n317_), .B2(new_n285_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n315_), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n318_), .A2(new_n319_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT101), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n324_));
  NAND2_X1  g123(.A1(new_n297_), .A2(new_n271_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n256_), .B1(G183gat), .B2(G190gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n254_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n261_), .A2(KEYINPUT24), .A3(new_n249_), .ZN(new_n328_));
  XOR2_X1   g127(.A(KEYINPUT25), .B(G183gat), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n264_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n260_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n328_), .A2(new_n331_), .A3(new_n256_), .A4(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n327_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n295_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT98), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n340_), .A2(KEYINPUT20), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n336_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT98), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AND4_X1   g143(.A1(new_n325_), .A2(new_n337_), .A3(new_n341_), .A4(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT20), .B1(new_n297_), .B2(new_n271_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT97), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n297_), .C2(new_n271_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n335_), .A2(new_n336_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n340_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n345_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT18), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  NOR2_X1   g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n357_), .ZN(new_n359_));
  AOI211_X1 g158(.A(new_n359_), .B(new_n345_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n324_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n353_), .A2(new_n357_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n348_), .A2(new_n340_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n325_), .A2(KEYINPUT20), .A3(new_n342_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n352_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n362_), .B(KEYINPUT27), .C1(new_n357_), .C2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n322_), .A2(new_n323_), .A3(new_n361_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n361_), .A2(new_n367_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT101), .B1(new_n369_), .B2(new_n321_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n283_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT99), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n234_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n245_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT33), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n244_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n239_), .A2(KEYINPUT33), .A3(new_n243_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n358_), .A2(new_n360_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n357_), .A2(KEYINPUT32), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n380_), .B2(new_n353_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n378_), .A2(new_n379_), .B1(new_n247_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n372_), .B1(new_n383_), .B2(new_n321_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n353_), .A2(new_n357_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n385_), .A2(new_n376_), .A3(new_n362_), .A4(new_n377_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n247_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n321_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT99), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n321_), .A2(new_n361_), .A3(new_n248_), .A4(new_n367_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n384_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n282_), .A2(KEYINPUT90), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n282_), .A2(KEYINPUT90), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n371_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G29gat), .B(G36gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G43gat), .B(G50gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT15), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G15gat), .B(G22gat), .ZN(new_n400_));
  INV_X1    g199(.A(G1gat), .ZN(new_n401_));
  INV_X1    g200(.A(G8gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT14), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT77), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n400_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n403_), .A2(new_n404_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G1gat), .B(G8gat), .ZN(new_n407_));
  OR3_X1    g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n399_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G229gat), .A2(G233gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n409_), .A3(new_n398_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n412_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n413_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n398_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G113gat), .B(G141gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G169gat), .B(G197gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  NAND3_X1  g220(.A1(new_n414_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT81), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI211_X1 g224(.A(KEYINPUT81), .B(new_n421_), .C1(new_n414_), .C2(new_n418_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT82), .Z(new_n428_));
  XNOR2_X1  g227(.A(G85gat), .B(G92gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT6), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(G99gat), .A3(G106gat), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n431_), .A2(new_n433_), .A3(KEYINPUT71), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT71), .B1(new_n431_), .B2(new_n433_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT68), .B1(G99gat), .B2(G106gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT7), .B1(new_n437_), .B2(KEYINPUT69), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT68), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n429_), .B1(new_n436_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT8), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT72), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n431_), .A2(new_n433_), .ZN(new_n448_));
  AOI211_X1 g247(.A(G99gat), .B(G106gat), .C1(new_n440_), .C2(KEYINPUT68), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n438_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT70), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n429_), .A2(KEYINPUT8), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT72), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n437_), .A2(KEYINPUT69), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n457_), .A2(new_n458_), .B1(new_n442_), .B2(new_n441_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n459_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n456_), .B(KEYINPUT8), .C1(new_n460_), .C2(new_n429_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n447_), .A2(new_n455_), .A3(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G64gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT73), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G71gat), .B(G78gat), .Z(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(KEYINPUT11), .B2(new_n463_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n466_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT9), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n429_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT10), .B(G99gat), .Z(new_n472_));
  INV_X1    g271(.A(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT66), .B(G92gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n470_), .A3(G85gat), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n471_), .A2(new_n474_), .A3(new_n448_), .A4(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n477_), .B(KEYINPUT67), .Z(new_n478_));
  AND3_X1   g277(.A1(new_n462_), .A2(new_n469_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n469_), .B1(new_n462_), .B2(new_n478_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT12), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G230gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n462_), .A2(new_n478_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n469_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT12), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(new_n484_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n462_), .A2(new_n469_), .A3(new_n478_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n484_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G120gat), .B(G148gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT5), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G176gat), .B(G204gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n490_), .A2(new_n494_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT74), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(KEYINPUT74), .A3(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n508_), .A2(KEYINPUT13), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(KEYINPUT13), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n395_), .A2(new_n428_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT34), .Z(new_n514_));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT75), .Z(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT76), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n485_), .B2(new_n399_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n398_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n485_), .B2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n514_), .A2(new_n515_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G134gat), .B(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n526_), .A2(KEYINPUT36), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(KEYINPUT36), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n523_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT37), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n410_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(new_n469_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G127gat), .B(G155gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G183gat), .B(G211gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT80), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT78), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n536_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n536_), .A2(new_n546_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n543_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n533_), .A2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n512_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(new_n401_), .A3(new_n247_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT38), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT102), .Z(new_n557_));
  INV_X1    g356(.A(new_n531_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n395_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n511_), .ZN(new_n560_));
  AND4_X1   g359(.A1(new_n550_), .A2(new_n559_), .A3(new_n427_), .A4(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n401_), .B1(new_n561_), .B2(new_n247_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n555_), .B2(new_n554_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n563_), .ZN(G1324gat));
  AOI21_X1  g363(.A(new_n402_), .B1(new_n561_), .B2(new_n369_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT39), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n553_), .A2(new_n402_), .A3(new_n369_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT40), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(KEYINPUT40), .A3(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(G1325gat));
  INV_X1    g372(.A(new_n394_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n278_), .B1(new_n561_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n553_), .A2(new_n278_), .A3(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(G1326gat));
  INV_X1    g378(.A(G22gat), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n561_), .B2(new_n321_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT42), .Z(new_n582_));
  NAND3_X1  g381(.A1(new_n553_), .A2(new_n580_), .A3(new_n321_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(G1327gat));
  NOR2_X1   g383(.A1(new_n531_), .A2(new_n550_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n512_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(G29gat), .B1(new_n586_), .B2(new_n247_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT104), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT43), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT43), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n531_), .B(KEYINPUT37), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n589_), .B(new_n590_), .C1(new_n395_), .C2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n390_), .B1(new_n388_), .B2(KEYINPUT99), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n383_), .A2(new_n372_), .A3(new_n321_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n394_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n371_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n597_), .A2(new_n588_), .A3(KEYINPUT43), .A4(new_n533_), .ZN(new_n598_));
  NOR4_X1   g397(.A1(new_n511_), .A2(new_n550_), .A3(new_n426_), .A4(new_n425_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n592_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT44), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT105), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(KEYINPUT105), .A3(new_n601_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n247_), .A2(G29gat), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n587_), .B1(new_n607_), .B2(new_n608_), .ZN(G1328gat));
  INV_X1    g408(.A(G36gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n607_), .B2(new_n369_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n586_), .A2(new_n610_), .A3(new_n369_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT45), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(G1329gat));
  INV_X1    g419(.A(new_n602_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n282_), .ZN(new_n622_));
  INV_X1    g421(.A(G43gat), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n600_), .A2(KEYINPUT105), .A3(new_n601_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT105), .B1(new_n600_), .B2(new_n601_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n621_), .B(new_n624_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT107), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n605_), .A2(new_n606_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT107), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n621_), .A4(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n586_), .A2(new_n574_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n623_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n628_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT47), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT47), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n628_), .A2(new_n631_), .A3(new_n636_), .A4(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1330gat));
  AOI21_X1  g437(.A(G50gat), .B1(new_n586_), .B2(new_n321_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n321_), .A2(G50gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n607_), .B2(new_n640_), .ZN(G1331gat));
  NAND2_X1  g440(.A1(new_n428_), .A2(new_n550_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n560_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n559_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G57gat), .B1(new_n645_), .B2(new_n248_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n395_), .A2(new_n427_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT108), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n552_), .A3(new_n511_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n248_), .A2(G57gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1332gat));
  INV_X1    g450(.A(G64gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n644_), .B2(new_n369_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT48), .Z(new_n654_));
  NAND2_X1  g453(.A1(new_n369_), .A2(new_n652_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n649_), .B2(new_n655_), .ZN(G1333gat));
  INV_X1    g455(.A(G71gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n644_), .B2(new_n574_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n574_), .A2(new_n657_), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n660_), .A2(new_n661_), .B1(new_n649_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT110), .ZN(G1334gat));
  INV_X1    g463(.A(G78gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n644_), .B2(new_n321_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT50), .Z(new_n667_));
  NAND2_X1  g466(.A1(new_n321_), .A2(new_n665_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n649_), .B2(new_n668_), .ZN(G1335gat));
  AND3_X1   g468(.A1(new_n648_), .A2(new_n511_), .A3(new_n585_), .ZN(new_n670_));
  INV_X1    g469(.A(G85gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n671_), .A3(new_n247_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n560_), .A2(new_n550_), .A3(new_n427_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n592_), .A2(new_n598_), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT111), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT112), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n676_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n248_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n672_), .B1(new_n679_), .B2(new_n671_), .ZN(G1336gat));
  AOI21_X1  g479(.A(G92gat), .B1(new_n670_), .B2(new_n369_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n677_), .A2(new_n678_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n369_), .A2(new_n475_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(G1337gat));
  NAND2_X1  g483(.A1(new_n675_), .A2(new_n574_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n282_), .A2(new_n472_), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n685_), .A2(G99gat), .B1(new_n670_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT51), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1338gat));
  OR2_X1    g488(.A1(new_n674_), .A2(new_n322_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(G106gat), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT52), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n322_), .A2(G106gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT113), .B1(new_n670_), .B2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n648_), .A2(new_n511_), .A3(new_n585_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT113), .ZN(new_n698_));
  INV_X1    g497(.A(new_n695_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n691_), .B(new_n694_), .C1(new_n696_), .C2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT53), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n670_), .A2(KEYINPUT113), .A3(new_n695_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT53), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n691_), .A4(new_n694_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n702_), .A2(new_n707_), .ZN(G1339gat));
  AOI211_X1 g507(.A(new_n248_), .B(new_n622_), .C1(new_n368_), .C2(new_n370_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT57), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n411_), .A2(new_n415_), .A3(new_n413_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n412_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n421_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n422_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n507_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n502_), .A2(new_n427_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT115), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n480_), .A2(KEYINPUT12), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n492_), .B2(KEYINPUT12), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT116), .B1(new_n720_), .B2(new_n484_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n481_), .A2(new_n489_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT116), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n493_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT55), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n490_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n481_), .A2(KEYINPUT55), .A3(new_n489_), .A4(new_n484_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n721_), .A2(new_n724_), .A3(new_n726_), .A4(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n728_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n499_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n718_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n499_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT56), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT117), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n728_), .A2(KEYINPUT56), .A3(new_n499_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n716_), .B1(new_n730_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n710_), .B1(new_n737_), .B2(new_n558_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n718_), .A2(new_n729_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n735_), .A2(new_n734_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n733_), .B2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT57), .B(new_n531_), .C1(new_n741_), .C2(new_n716_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n735_), .A2(KEYINPUT118), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT118), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n728_), .A2(new_n745_), .A3(KEYINPUT56), .A4(new_n499_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n744_), .A2(new_n746_), .A3(new_n733_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n715_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n502_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT58), .B1(new_n747_), .B2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT119), .B1(new_n751_), .B2(new_n591_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT119), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT56), .B1(new_n728_), .B2(new_n499_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(KEYINPUT118), .B2(new_n735_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n749_), .B1(new_n755_), .B2(new_n746_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n753_), .B(new_n533_), .C1(new_n756_), .C2(KEYINPUT58), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(KEYINPUT58), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n743_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n752_), .A2(new_n757_), .A3(KEYINPUT120), .A4(new_n758_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n550_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n533_), .A2(new_n642_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n560_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n765_), .B(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n709_), .B1(new_n763_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(G113gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n427_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT59), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n709_), .A2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n738_), .A2(new_n742_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n759_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n551_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n765_), .B(new_n766_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n428_), .B(new_n779_), .C1(new_n769_), .C2(KEYINPUT59), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n772_), .B1(new_n780_), .B2(new_n771_), .ZN(G1340gat));
  INV_X1    g580(.A(KEYINPUT121), .ZN(new_n782_));
  INV_X1    g581(.A(G120gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n779_), .B1(new_n769_), .B2(KEYINPUT59), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n511_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT60), .ZN(new_n786_));
  AOI21_X1  g585(.A(G120gat), .B1(new_n511_), .B2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n783_), .A2(KEYINPUT60), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n769_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n782_), .B1(new_n785_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n789_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n560_), .B(new_n779_), .C1(new_n769_), .C2(KEYINPUT59), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n791_), .B(KEYINPUT121), .C1(new_n792_), .C2(new_n783_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1341gat));
  INV_X1    g593(.A(G127gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n770_), .A2(new_n795_), .A3(new_n550_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n784_), .A2(new_n550_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n795_), .ZN(G1342gat));
  INV_X1    g597(.A(G134gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n770_), .A2(new_n799_), .A3(new_n558_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n784_), .A2(new_n533_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n799_), .ZN(G1343gat));
  OR2_X1    g601(.A1(new_n763_), .A2(new_n768_), .ZN(new_n803_));
  NOR4_X1   g602(.A1(new_n574_), .A2(new_n369_), .A3(new_n322_), .A4(new_n248_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n427_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n511_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g608(.A1(new_n803_), .A2(new_n804_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n551_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT61), .B(G155gat), .Z(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(G1346gat));
  OAI211_X1 g612(.A(new_n533_), .B(new_n804_), .C1(new_n763_), .C2(new_n768_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G162gat), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n531_), .A2(G162gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n810_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT122), .ZN(G1347gat));
  AOI21_X1  g617(.A(new_n550_), .B1(new_n775_), .B2(new_n759_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n768_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n369_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n821_), .A2(new_n394_), .A3(new_n247_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n322_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT123), .B1(new_n820_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n777_), .A2(new_n778_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT123), .ZN(new_n826_));
  INV_X1    g625(.A(new_n823_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n251_), .A3(new_n427_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n825_), .A2(new_n427_), .A3(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G169gat), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n832_), .A2(KEYINPUT62), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(KEYINPUT62), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n830_), .B1(new_n833_), .B2(new_n834_), .ZN(G1348gat));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  INV_X1    g635(.A(new_n829_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n836_), .B(new_n252_), .C1(new_n837_), .C2(new_n560_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n560_), .B1(new_n824_), .B2(new_n828_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT124), .B1(new_n839_), .B2(G176gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n763_), .A2(new_n768_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT125), .B1(new_n841_), .B2(new_n321_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n843_), .B(new_n322_), .C1(new_n763_), .C2(new_n768_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n842_), .A2(new_n822_), .A3(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n560_), .A2(new_n252_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n838_), .A2(new_n840_), .B1(new_n845_), .B2(new_n846_), .ZN(G1349gat));
  NAND4_X1  g646(.A1(new_n842_), .A2(new_n550_), .A3(new_n822_), .A4(new_n844_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n257_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n551_), .A2(new_n330_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n848_), .A2(new_n849_), .B1(new_n829_), .B2(new_n850_), .ZN(G1350gat));
  OAI21_X1  g650(.A(G190gat), .B1(new_n837_), .B2(new_n591_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n829_), .A2(new_n558_), .A3(new_n264_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1351gat));
  NAND3_X1  g653(.A1(new_n394_), .A2(new_n321_), .A3(new_n248_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT126), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n841_), .A2(new_n821_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n427_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n511_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n856_), .A2(new_n821_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n803_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n864_), .B2(new_n551_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT127), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT127), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n867_), .B(new_n862_), .C1(new_n864_), .C2(new_n551_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n864_), .A2(new_n551_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT63), .B(G211gat), .Z(new_n870_));
  AOI22_X1  g669(.A1(new_n866_), .A2(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1354gat));
  OAI21_X1  g670(.A(G218gat), .B1(new_n864_), .B2(new_n591_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n531_), .A2(G218gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n864_), .B2(new_n873_), .ZN(G1355gat));
endmodule


