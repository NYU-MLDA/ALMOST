//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT13), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT10), .B(G99gat), .Z(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT65), .Z(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n212_), .A2(KEYINPUT9), .A3(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n217_), .B(KEYINPUT6), .Z(new_n218_));
  NOR3_X1   g017(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n208_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT67), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n222_), .B(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(new_n218_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n230_), .A3(new_n215_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n226_), .B2(new_n215_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n220_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT69), .ZN(new_n237_));
  XOR2_X1   g036(.A(G71gat), .B(G78gat), .Z(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(KEYINPUT11), .B2(new_n235_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n234_), .A2(new_n241_), .A3(KEYINPUT12), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n226_), .A2(new_n215_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n229_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n244_), .A2(new_n231_), .B1(new_n219_), .B2(new_n210_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n240_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT64), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n234_), .A2(new_n241_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT12), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT70), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n244_), .A2(new_n231_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n240_), .B1(new_n254_), .B2(new_n220_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n255_), .A2(new_n256_), .A3(KEYINPUT12), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n248_), .B(new_n250_), .C1(new_n253_), .C2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n255_), .B2(KEYINPUT12), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n251_), .A2(KEYINPUT70), .A3(new_n252_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n247_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(KEYINPUT71), .A3(new_n250_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n246_), .A2(new_n251_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n250_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G120gat), .B(G148gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT5), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G176gat), .B(G204gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT72), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n268_), .A3(new_n274_), .ZN(new_n277_));
  AOI211_X1 g076(.A(new_n205_), .B(new_n206_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n276_), .A2(KEYINPUT73), .A3(KEYINPUT13), .A4(new_n277_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n202_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n277_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n205_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n206_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(KEYINPUT74), .A3(new_n279_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G22gat), .B(G50gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT85), .B1(new_n301_), .B2(KEYINPUT3), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n300_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n295_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n293_), .B1(KEYINPUT1), .B2(new_n291_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n291_), .A2(KEYINPUT1), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n301_), .A3(new_n296_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT87), .B1(new_n311_), .B2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n298_), .A2(new_n299_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n306_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n304_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n308_), .B(KEYINPUT86), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n294_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n315_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n290_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(new_n329_), .A3(new_n289_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT92), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT92), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G211gat), .B(G218gat), .Z(new_n339_));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n340_));
  AND2_X1   g139(.A1(G197gat), .A2(G204gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G197gat), .A2(G204gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G197gat), .ZN(new_n344_));
  INV_X1    g143(.A(G204gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(KEYINPUT90), .A3(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n339_), .A2(new_n343_), .A3(new_n348_), .A4(KEYINPUT21), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT21), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n346_), .A2(KEYINPUT21), .A3(new_n347_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT88), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n346_), .A2(KEYINPUT88), .A3(KEYINPUT21), .A4(new_n347_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n349_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G228gat), .ZN(new_n361_));
  INV_X1    g160(.A(G233gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n317_), .A2(new_n325_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(KEYINPUT29), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n311_), .A2(new_n316_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n360_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n361_), .A2(new_n362_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(G78gat), .B1(new_n365_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G78gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n369_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n326_), .A2(new_n328_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n372_), .B(new_n373_), .C1(new_n374_), .C2(new_n363_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n208_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n208_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n336_), .B(new_n338_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n380_), .A2(KEYINPUT92), .A3(new_n335_), .A4(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G127gat), .B(G134gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G113gat), .B(G120gat), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n390_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n391_), .A2(KEYINPUT84), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT84), .B1(new_n391_), .B2(new_n392_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n317_), .A2(new_n325_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n366_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT4), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n388_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n396_), .A2(new_n388_), .A3(new_n398_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT98), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n396_), .A2(KEYINPUT98), .A3(new_n388_), .A4(new_n398_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n387_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n388_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n402_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n401_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n387_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n406_), .A4(new_n407_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G183gat), .ZN(new_n422_));
  INV_X1    g221(.A(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G169gat), .ZN(new_n425_));
  OR3_X1    g224(.A1(new_n425_), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n421_), .A2(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT25), .B(G183gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G190gat), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT83), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT83), .B1(new_n429_), .B2(new_n430_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n419_), .A2(new_n434_), .A3(new_n420_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G169gat), .A2(G176gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n428_), .B1(new_n433_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(G15gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT30), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n441_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(new_n395_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G43gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT31), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n447_), .B(new_n451_), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n417_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n420_), .ZN(new_n454_));
  INV_X1    g253(.A(G176gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n425_), .A2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n454_), .B(new_n418_), .C1(new_n456_), .C2(KEYINPUT24), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n422_), .A2(KEYINPUT25), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G183gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n423_), .A2(KEYINPUT26), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT26), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G190gat), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n458_), .A2(new_n460_), .A3(new_n461_), .A4(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n439_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n457_), .B1(new_n465_), .B2(KEYINPUT94), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n429_), .A2(new_n430_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT94), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n428_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n349_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n351_), .B(KEYINPUT89), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT95), .B1(new_n470_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n441_), .B2(new_n474_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n428_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n435_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n465_), .A2(KEYINPUT94), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n360_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n477_), .A3(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G226gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT96), .ZN(new_n490_));
  XOR2_X1   g289(.A(G8gat), .B(G36gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT20), .B1(new_n481_), .B2(new_n360_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n441_), .A2(new_n474_), .ZN(new_n498_));
  OR3_X1    g297(.A1(new_n497_), .A2(new_n498_), .A3(new_n488_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n484_), .A2(new_n500_), .A3(new_n488_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n490_), .A2(new_n496_), .A3(new_n499_), .A4(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT27), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n488_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n503_), .B1(new_n505_), .B2(new_n495_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n499_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n500_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n495_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n502_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT102), .B1(new_n511_), .B2(new_n503_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT102), .ZN(new_n513_));
  AOI211_X1 g312(.A(new_n513_), .B(KEYINPUT27), .C1(new_n510_), .C2(new_n502_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n507_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT103), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT103), .B(new_n507_), .C1(new_n512_), .C2(new_n514_), .ZN(new_n518_));
  AOI211_X1 g317(.A(new_n383_), .B(new_n453_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n510_), .A2(new_n502_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n513_), .B1(new_n520_), .B2(KEYINPUT27), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n511_), .A2(KEYINPUT102), .A3(new_n503_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n523_), .A2(new_n383_), .A3(new_n417_), .A4(new_n507_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n388_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n387_), .C1(new_n388_), .C2(new_n399_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT33), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n387_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n413_), .A2(new_n406_), .A3(new_n407_), .A4(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n510_), .A2(new_n527_), .A3(new_n502_), .A4(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n403_), .A2(new_n408_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT33), .B1(new_n532_), .B2(new_n414_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n525_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n387_), .B1(new_n399_), .B2(new_n388_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n400_), .A2(new_n402_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n388_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n532_), .B2(new_n529_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n415_), .A2(new_n528_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n520_), .A2(KEYINPUT99), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n495_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n505_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT101), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n542_), .B(KEYINPUT100), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n490_), .A2(new_n545_), .A3(new_n499_), .A4(new_n501_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT101), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n505_), .A2(new_n547_), .A3(new_n542_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n544_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n416_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n534_), .A2(new_n540_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n382_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n452_), .B1(new_n524_), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n519_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT80), .B(G8gat), .Z(new_n555_));
  INV_X1    g354(.A(G1gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT79), .B(G15gat), .ZN(new_n558_));
  INV_X1    g357(.A(G22gat), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n559_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G1gat), .B(G8gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(G29gat), .B(G36gat), .Z(new_n568_));
  XOR2_X1   g367(.A(G43gat), .B(G50gat), .Z(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n567_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n570_), .B(KEYINPUT15), .Z(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n570_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n567_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n577_), .A3(new_n572_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n573_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n554_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT77), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n254_), .A2(new_n570_), .A3(new_n220_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n245_), .B2(new_n574_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT35), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(KEYINPUT76), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(KEYINPUT35), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n590_), .B2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT76), .B1(new_n590_), .B2(new_n593_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n588_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT75), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(G134gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G162gat), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n602_), .A2(new_n603_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  OAI221_X1 g407(.A(new_n588_), .B1(new_n606_), .B2(new_n604_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT78), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT37), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT78), .B(new_n613_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n567_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n240_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT17), .ZN(new_n620_));
  XOR2_X1   g419(.A(G127gat), .B(G155gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n619_), .A2(new_n620_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT82), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n625_), .B(KEYINPUT17), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n619_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n615_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n288_), .A2(new_n587_), .A3(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT104), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(KEYINPUT104), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n633_), .A2(new_n556_), .A3(new_n416_), .A4(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n637_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n554_), .A2(new_n610_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n285_), .A2(new_n279_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n641_), .A2(new_n586_), .A3(new_n630_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n417_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n638_), .A2(new_n639_), .A3(new_n644_), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n517_), .A2(new_n518_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(new_n555_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n633_), .A2(new_n634_), .A3(new_n648_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n643_), .A2(KEYINPUT106), .A3(new_n646_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT106), .B1(new_n643_), .B2(new_n646_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(G8gat), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n650_), .A2(new_n654_), .A3(G8gat), .A4(new_n651_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n649_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n656_), .B(new_n658_), .ZN(G1325gat));
  INV_X1    g458(.A(new_n452_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G15gat), .B1(new_n643_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n632_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n443_), .A3(new_n452_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n664_), .A3(new_n666_), .ZN(G1326gat));
  OAI21_X1  g466(.A(G22gat), .B1(new_n643_), .B2(new_n382_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT42), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n559_), .A3(new_n383_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1327gat));
  NOR2_X1   g470(.A1(new_n278_), .A2(new_n280_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n630_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n610_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n587_), .A2(new_n672_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT111), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT111), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n587_), .A2(new_n672_), .A3(new_n678_), .A4(new_n675_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n416_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n586_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n672_), .A2(new_n682_), .A3(new_n630_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n684_));
  NOR2_X1   g483(.A1(new_n612_), .A2(new_n614_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n554_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n687_), .B(new_n615_), .C1(new_n519_), .C2(new_n553_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n683_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT110), .B1(new_n689_), .B2(KEYINPUT44), .ZN(new_n690_));
  INV_X1    g489(.A(new_n453_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n646_), .A2(new_n382_), .A3(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n538_), .A2(new_n502_), .A3(new_n510_), .A4(new_n539_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n693_), .A2(new_n525_), .B1(new_n416_), .B2(new_n549_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n383_), .B1(new_n694_), .B2(new_n540_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n379_), .A2(new_n381_), .A3(new_n417_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n515_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n660_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n685_), .B1(new_n692_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n684_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n688_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n641_), .A2(new_n586_), .A3(new_n673_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n690_), .A2(new_n706_), .B1(KEYINPUT44), .B2(new_n689_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n416_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n681_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n677_), .A2(new_n710_), .A3(new_n647_), .A4(new_n679_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n701_), .A2(KEYINPUT44), .A3(new_n702_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n647_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n690_), .B2(new_n706_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n710_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n646_), .B1(new_n689_), .B2(KEYINPUT44), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n704_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n701_), .C2(new_n702_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT112), .B1(new_n722_), .B2(G36gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n713_), .B1(new_n718_), .B2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI221_X1 g525(.A(new_n713_), .B1(KEYINPUT114), .B2(KEYINPUT46), .C1(new_n718_), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  NAND3_X1  g527(.A1(new_n707_), .A2(G43gat), .A3(new_n452_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n680_), .A2(new_n452_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n449_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n680_), .B2(new_n383_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n383_), .A2(G50gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n707_), .B2(new_n735_), .ZN(G1331gat));
  NAND4_X1  g535(.A1(new_n640_), .A2(new_n287_), .A3(new_n586_), .A4(new_n673_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n417_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n554_), .A2(new_n682_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n739_), .A2(new_n641_), .A3(new_n631_), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n416_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n744_), .A3(new_n647_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G64gat), .B1(new_n737_), .B2(new_n646_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT48), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT48), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n740_), .A2(new_n750_), .A3(new_n452_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G71gat), .B1(new_n737_), .B2(new_n660_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(KEYINPUT116), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n751_), .B1(new_n756_), .B2(new_n757_), .ZN(G1334gat));
  NAND3_X1  g557(.A1(new_n740_), .A2(new_n372_), .A3(new_n383_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G78gat), .B1(new_n737_), .B2(new_n382_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT50), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT50), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1335gat));
  NAND3_X1  g562(.A1(new_n739_), .A2(new_n287_), .A3(new_n675_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n416_), .ZN(new_n766_));
  AND4_X1   g565(.A1(new_n586_), .A2(new_n701_), .A3(new_n641_), .A4(new_n630_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n417_), .A2(new_n212_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(G1336gat));
  NAND3_X1  g568(.A1(new_n765_), .A2(new_n213_), .A3(new_n647_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n767_), .A2(new_n647_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n213_), .ZN(G1337gat));
  NAND2_X1  g571(.A1(new_n452_), .A2(new_n207_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n764_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT117), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n221_), .B1(new_n767_), .B2(new_n452_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g577(.A1(new_n765_), .A2(new_n208_), .A3(new_n383_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n767_), .A2(new_n383_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(G106gat), .ZN(new_n782_));
  AOI211_X1 g581(.A(KEYINPUT52), .B(new_n208_), .C1(new_n767_), .C2(new_n383_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT121), .ZN(new_n787_));
  INV_X1    g586(.A(new_n273_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n265_), .A2(new_n268_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n682_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n248_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT119), .A3(new_n267_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n263_), .B2(new_n250_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n267_), .B(new_n247_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n792_), .A2(new_n794_), .B1(new_n795_), .B2(KEYINPUT55), .ZN(new_n796_));
  XOR2_X1   g595(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n797_));
  NAND3_X1  g596(.A1(new_n260_), .A2(new_n264_), .A3(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n796_), .A2(KEYINPUT120), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT120), .B1(new_n796_), .B2(new_n798_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n273_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n792_), .A2(new_n794_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n795_), .A2(KEYINPUT55), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n798_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n796_), .A2(KEYINPUT120), .A3(new_n798_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n273_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n790_), .B1(new_n803_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n572_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n575_), .A2(new_n577_), .A3(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n814_), .B(new_n583_), .C1(new_n571_), .C2(new_n813_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n585_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n282_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n674_), .B(new_n787_), .C1(new_n812_), .C2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n789_), .A2(new_n816_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n273_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n802_), .B(new_n788_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT58), .B(new_n820_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n615_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n803_), .A2(new_n811_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT58), .B1(new_n825_), .B2(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n819_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n821_), .A2(new_n822_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n817_), .B1(new_n828_), .B2(new_n790_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n787_), .B1(new_n829_), .B2(new_n674_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n630_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n685_), .A2(new_n586_), .A3(new_n673_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n641_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT54), .Z(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n646_), .A2(new_n416_), .A3(new_n382_), .A4(new_n452_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT122), .Z(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(G113gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n682_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n838_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n835_), .A2(KEYINPUT59), .A3(new_n837_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n586_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n845_), .B2(new_n840_), .ZN(G1340gat));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n672_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n839_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n288_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n847_), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n839_), .B2(new_n673_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n843_), .A2(new_n844_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n630_), .A2(KEYINPUT123), .ZN(new_n854_));
  MUX2_X1   g653(.A(KEYINPUT123), .B(new_n854_), .S(G127gat), .Z(new_n855_));
  AOI21_X1  g654(.A(new_n852_), .B1(new_n853_), .B2(new_n855_), .ZN(G1342gat));
  INV_X1    g655(.A(G134gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n839_), .A2(new_n857_), .A3(new_n610_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n685_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n857_), .ZN(G1343gat));
  NOR3_X1   g659(.A1(new_n647_), .A2(new_n417_), .A3(new_n382_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n452_), .B(new_n862_), .C1(new_n831_), .C2(new_n834_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n682_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n287_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n863_), .B2(new_n673_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n835_), .A2(new_n660_), .A3(new_n673_), .A4(new_n861_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(KEYINPUT124), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n869_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n863_), .A2(new_n870_), .A3(new_n673_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(KEYINPUT124), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n868_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(new_n877_), .ZN(G1346gat));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n863_), .A2(new_n879_), .A3(new_n610_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n835_), .A2(new_n660_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n881_), .A2(new_n685_), .A3(new_n862_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n882_), .B2(new_n879_), .ZN(G1347gat));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n383_), .A2(new_n453_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n647_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n682_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n888_), .B2(G169gat), .ZN(new_n889_));
  AOI211_X1 g688(.A(KEYINPUT62), .B(new_n425_), .C1(new_n887_), .C2(new_n682_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n887_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT22), .B(G169gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n682_), .A2(new_n892_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT125), .Z(new_n894_));
  OAI22_X1  g693(.A1(new_n889_), .A2(new_n890_), .B1(new_n891_), .B2(new_n894_), .ZN(G1348gat));
  OAI21_X1  g694(.A(G176gat), .B1(new_n891_), .B2(new_n288_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n887_), .A2(new_n455_), .A3(new_n641_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1349gat));
  AOI21_X1  g697(.A(G183gat), .B1(new_n887_), .B2(new_n673_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n887_), .A2(new_n673_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n900_), .B(new_n901_), .C1(new_n429_), .C2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n429_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT126), .B1(new_n904_), .B2(new_n899_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n891_), .B2(new_n685_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n887_), .A2(new_n430_), .A3(new_n610_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1351gat));
  NOR2_X1   g708(.A1(new_n646_), .A2(new_n696_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n881_), .A2(new_n586_), .A3(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n344_), .ZN(G1352gat));
  NOR3_X1   g712(.A1(new_n881_), .A2(new_n288_), .A3(new_n911_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n345_), .ZN(G1353gat));
  AOI21_X1  g714(.A(new_n630_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n835_), .A2(new_n660_), .A3(new_n910_), .A4(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(KEYINPUT127), .B2(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(KEYINPUT127), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n917_), .B2(new_n920_), .ZN(G1354gat));
  OR4_X1    g720(.A1(G218gat), .A2(new_n881_), .A3(new_n674_), .A4(new_n911_), .ZN(new_n922_));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n881_), .A2(new_n685_), .A3(new_n911_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1355gat));
endmodule


