//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  XOR2_X1   g000(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT13), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT67), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(KEYINPUT67), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G230gat), .A2(G233gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT6), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  OR3_X1    g011(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G85gat), .B(G92gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n215_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT64), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n214_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT8), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G85gat), .ZN(new_n226_));
  INV_X1    g025(.A(G92gat), .ZN(new_n227_));
  OR3_X1    g026(.A1(new_n226_), .A2(new_n227_), .A3(KEYINPUT9), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n222_), .A2(new_n225_), .A3(new_n211_), .A4(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n221_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n232_));
  XOR2_X1   g031(.A(G71gat), .B(G78gat), .Z(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n233_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n230_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n221_), .A2(new_n229_), .A3(new_n237_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n239_), .A2(new_n240_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n209_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(KEYINPUT12), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n238_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n234_), .B(KEYINPUT12), .C1(new_n235_), .C2(new_n236_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n229_), .B1(new_n221_), .B2(KEYINPUT66), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n248_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n246_), .A2(new_n254_), .A3(new_n208_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G120gat), .B(G148gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT5), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G176gat), .B(G204gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n244_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n244_), .B2(new_n255_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n205_), .B(new_n207_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT13), .A4(new_n261_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G22gat), .ZN(new_n270_));
  INV_X1    g069(.A(G1gat), .ZN(new_n271_));
  INV_X1    g070(.A(G8gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT14), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G8gat), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n275_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G43gat), .B(G50gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(G29gat), .B(G36gat), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(KEYINPUT15), .Z(new_n285_));
  AOI21_X1  g084(.A(new_n284_), .B1(new_n285_), .B2(new_n278_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G229gat), .A2(G233gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n278_), .B(new_n283_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(new_n287_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G113gat), .B(G141gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(G169gat), .B(G197gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n292_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n269_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G134gat), .Z(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(new_n299_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT74), .B1(new_n302_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n301_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n299_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT31), .Z(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(G183gat), .B2(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n315_));
  OAI22_X1  g114(.A1(new_n313_), .A2(new_n315_), .B1(G183gat), .B2(G190gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT73), .B(G176gat), .ZN(new_n317_));
  INV_X1    g116(.A(G169gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT22), .B1(new_n318_), .B2(KEYINPUT72), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT22), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(G169gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(G169gat), .B2(G176gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n326_), .A2(new_n327_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n328_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n333_), .B(new_n334_), .C1(new_n313_), .C2(new_n315_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n312_), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n337_), .A2(new_n338_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(new_n333_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n325_), .B1(new_n336_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT30), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G71gat), .B(G99gat), .ZN(new_n343_));
  INV_X1    g142(.A(G43gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(G15gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n345_), .B(new_n348_), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n342_), .B(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n311_), .B1(new_n351_), .B2(KEYINPUT75), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n342_), .B(new_n349_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n354_), .A3(new_n311_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT0), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G57gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(G57gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n226_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n363_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G85gat), .A3(new_n361_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT2), .ZN(new_n368_));
  INV_X1    g167(.A(G141gat), .ZN(new_n369_));
  INV_X1    g168(.A(G148gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .A4(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT76), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n381_), .A3(new_n378_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n376_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G141gat), .B(G148gat), .Z(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(KEYINPUT1), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n377_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n378_), .A2(KEYINPUT1), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n384_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n383_), .A2(new_n308_), .A3(new_n306_), .A4(new_n388_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(KEYINPUT4), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n389_), .A2(new_n305_), .A3(new_n395_), .A4(new_n309_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n390_), .A2(new_n393_), .A3(new_n391_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n367_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n398_), .A3(new_n367_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n358_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n389_), .A2(KEYINPUT29), .ZN(new_n404_));
  INV_X1    g203(.A(G197gat), .ZN(new_n405_));
  INV_X1    g204(.A(G204gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(KEYINPUT21), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n407_), .A2(KEYINPUT82), .A3(KEYINPUT21), .A4(new_n408_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT21), .ZN(new_n413_));
  INV_X1    g212(.A(new_n408_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G197gat), .A2(G204gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G218gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G211gat), .ZN(new_n418_));
  INV_X1    g217(.A(G211gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G218gat), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n411_), .A2(new_n412_), .A3(new_n416_), .A4(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n409_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n418_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n423_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n404_), .A2(KEYINPUT81), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G228gat), .A2(G233gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n430_), .B(KEYINPUT80), .Z(new_n431_));
  XNOR2_X1  g230(.A(new_n429_), .B(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT77), .B(KEYINPUT28), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n389_), .A2(KEYINPUT29), .A3(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n435_), .B1(new_n389_), .B2(KEYINPUT29), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT78), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT79), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n436_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT84), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n443_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n445_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n433_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n444_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n441_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n445_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n443_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n432_), .A3(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT19), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT22), .B(G169gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n317_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n316_), .A2(new_n324_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G183gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT25), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT25), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(G183gat), .ZN(new_n466_));
  INV_X1    g265(.A(G190gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT26), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT26), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(G190gat), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n464_), .A2(new_n466_), .A3(new_n468_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n329_), .A2(new_n331_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n339_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n462_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT20), .B1(new_n428_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n334_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT71), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(new_n335_), .A3(new_n332_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n478_), .A2(new_n325_), .B1(new_n422_), .B2(new_n427_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n459_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n339_), .A2(new_n471_), .A3(new_n472_), .A4(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n462_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n332_), .B2(new_n339_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n428_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n478_), .A2(new_n325_), .A3(new_n422_), .A4(new_n427_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT20), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n480_), .B1(new_n459_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G8gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT18), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G64gat), .B(G92gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT27), .ZN(new_n494_));
  INV_X1    g293(.A(new_n492_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n487_), .A2(new_n459_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n487_), .A2(KEYINPUT86), .A3(new_n459_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n473_), .A2(KEYINPUT85), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(new_n482_), .A3(new_n462_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n502_), .B2(new_n428_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n422_), .A2(new_n427_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n462_), .A2(new_n482_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT87), .A4(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n458_), .A2(KEYINPUT20), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n341_), .B2(new_n428_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT88), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n503_), .A2(new_n506_), .A3(new_n508_), .A4(KEYINPUT88), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n498_), .A2(new_n499_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n494_), .B1(new_n495_), .B2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n511_), .A2(new_n512_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n487_), .A2(KEYINPUT86), .A3(new_n459_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT86), .B1(new_n487_), .B2(new_n459_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n492_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n498_), .A2(new_n499_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n511_), .A2(new_n512_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n495_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT27), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n514_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n403_), .A2(new_n456_), .A3(new_n525_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n520_), .A2(new_n521_), .A3(new_n495_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n495_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n402_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n522_), .A2(KEYINPUT27), .A3(new_n493_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT89), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n529_), .A2(new_n530_), .A3(new_n534_), .A4(new_n531_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT33), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n401_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n397_), .A2(KEYINPUT33), .A3(new_n398_), .A4(new_n367_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n392_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n390_), .A2(new_n394_), .A3(new_n391_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n539_), .A2(new_n366_), .A3(new_n364_), .A4(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n527_), .A2(new_n528_), .A3(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n495_), .A2(KEYINPUT32), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n488_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n401_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n545_), .B1(new_n546_), .B2(new_n399_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n544_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n547_), .B1(new_n513_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n456_), .B1(new_n543_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n533_), .A2(new_n535_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n526_), .B1(new_n551_), .B2(new_n358_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n298_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G190gat), .B(G218gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT36), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n562_));
  INV_X1    g361(.A(new_n283_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n230_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n285_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n557_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n565_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n566_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n556_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(KEYINPUT36), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT69), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n278_), .B(new_n581_), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n237_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n583_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(KEYINPUT70), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT70), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n583_), .A2(new_n589_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n580_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n553_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT90), .Z(new_n598_));
  INV_X1    g397(.A(new_n402_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(G1gat), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n203_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT95), .Z(new_n602_));
  NOR2_X1   g401(.A1(new_n298_), .A2(new_n595_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n569_), .A2(new_n576_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n552_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT93), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n599_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT94), .Z(new_n610_));
  NAND3_X1  g409(.A1(new_n598_), .A2(new_n600_), .A3(new_n203_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT92), .Z(new_n612_));
  NAND3_X1  g411(.A1(new_n602_), .A2(new_n610_), .A3(new_n612_), .ZN(G1324gat));
  INV_X1    g412(.A(new_n525_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n598_), .A2(new_n272_), .A3(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n607_), .B2(new_n525_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT39), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g418(.A(G15gat), .B1(new_n608_), .B2(new_n358_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT41), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT41), .ZN(new_n622_));
  INV_X1    g421(.A(new_n358_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n598_), .A2(new_n347_), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n621_), .A2(new_n622_), .A3(new_n624_), .ZN(G1326gat));
  XNOR2_X1  g424(.A(new_n456_), .B(KEYINPUT96), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n608_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G22gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT97), .B(KEYINPUT42), .Z(new_n629_));
  OR3_X1    g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n626_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n598_), .A2(new_n628_), .A3(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT98), .ZN(G1327gat));
  INV_X1    g434(.A(new_n595_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n604_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n553_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n639_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n642_), .A2(G29gat), .A3(new_n599_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n578_), .B(KEYINPUT37), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n550_), .A2(new_n535_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n534_), .B1(new_n525_), .B2(new_n530_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n358_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n526_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n644_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NOR4_X1   g453(.A1(new_n552_), .A2(KEYINPUT99), .A3(KEYINPUT43), .A4(new_n645_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n298_), .A2(new_n636_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n657_), .A2(KEYINPUT44), .A3(new_n658_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n402_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n663_), .A2(new_n664_), .A3(G29gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n663_), .B2(G29gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n643_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT103), .B(new_n643_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1328gat));
  AND2_X1   g470(.A1(new_n661_), .A2(new_n662_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n614_), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(KEYINPUT104), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n640_), .A2(new_n674_), .A3(new_n614_), .A4(new_n641_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT104), .B1(new_n678_), .B2(KEYINPUT45), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n679_), .B1(KEYINPUT45), .B2(new_n678_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n676_), .A2(new_n677_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n677_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1329gat));
  NAND3_X1  g482(.A1(new_n672_), .A2(G43gat), .A3(new_n623_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n344_), .B1(new_n642_), .B2(new_n358_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g486(.A1(new_n642_), .A2(new_n626_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(G50gat), .ZN(new_n689_));
  INV_X1    g488(.A(new_n456_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n661_), .A2(G50gat), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n662_), .B2(new_n691_), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n269_), .A2(new_n297_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n552_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n645_), .A2(new_n636_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n402_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n269_), .A2(new_n595_), .A3(new_n297_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n606_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n599_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n702_), .ZN(G1332gat));
  OAI21_X1  g502(.A(G64gat), .B1(new_n701_), .B2(new_n525_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT48), .ZN(new_n705_));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n706_), .A3(new_n614_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n697_), .A2(new_n709_), .A3(new_n623_), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT105), .B(KEYINPUT49), .Z(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n701_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n623_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n714_), .B2(G71gat), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n709_), .B(new_n711_), .C1(new_n713_), .C2(new_n623_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n710_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT106), .Z(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n701_), .B2(new_n626_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n697_), .A2(new_n721_), .A3(new_n632_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT107), .Z(G1335gat));
  AOI21_X1  g523(.A(new_n655_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n693_), .A2(new_n595_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n599_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n693_), .A2(new_n694_), .A3(new_n637_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n226_), .A3(new_n402_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1336gat));
  OAI21_X1  g533(.A(G92gat), .B1(new_n729_), .B2(new_n525_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n227_), .A3(new_n614_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1337gat));
  AND2_X1   g536(.A1(new_n623_), .A2(new_n223_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT109), .B1(new_n732_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n729_), .A2(new_n358_), .ZN(new_n740_));
  INV_X1    g539(.A(G99gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT51), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n739_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1338gat));
  INV_X1    g545(.A(new_n726_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n552_), .A2(KEYINPUT43), .A3(new_n645_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n552_), .B2(new_n645_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n644_), .B2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n690_), .B(new_n747_), .C1(new_n750_), .C2(new_n655_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT110), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n657_), .A2(new_n754_), .A3(new_n690_), .A4(new_n747_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .A4(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT111), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n725_), .A2(new_n456_), .A3(new_n726_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n224_), .B1(new_n758_), .B2(new_n754_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n753_), .A4(new_n752_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n755_), .A2(G106gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n754_), .B1(new_n727_), .B2(new_n690_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT52), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n757_), .A2(new_n761_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n732_), .A2(new_n224_), .A3(new_n690_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT53), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n765_), .A2(new_n769_), .A3(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1339gat));
  NOR3_X1   g570(.A1(new_n614_), .A2(new_n599_), .A3(new_n358_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n262_), .A2(new_n296_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n255_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n246_), .A2(new_n254_), .A3(KEYINPUT55), .A4(new_n208_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n246_), .A2(new_n254_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n209_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n259_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n259_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n773_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n295_), .B1(new_n290_), .B2(new_n287_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n286_), .A2(new_n288_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n295_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n783_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n789_), .A2(new_n790_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n796_), .A2(KEYINPUT116), .A3(new_n793_), .A4(new_n791_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n263_), .B2(new_n262_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n782_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT117), .B1(new_n800_), .B2(new_n604_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n262_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n803_), .B(KEYINPUT58), .C1(new_n780_), .C2(new_n781_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n580_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n801_), .A2(new_n802_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n605_), .B1(new_n782_), .B2(new_n799_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT57), .B1(new_n810_), .B2(KEYINPUT117), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n636_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n264_), .A2(new_n267_), .A3(new_n296_), .ZN(new_n813_));
  OR4_X1    g612(.A1(KEYINPUT112), .A2(new_n696_), .A3(new_n813_), .A4(KEYINPUT54), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n596_), .A2(new_n269_), .A3(new_n815_), .A4(new_n296_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT112), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n696_), .B2(new_n813_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT113), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(KEYINPUT54), .C1(new_n696_), .C2(new_n813_), .ZN(new_n821_));
  AND4_X1   g620(.A1(new_n814_), .A2(new_n817_), .A3(new_n819_), .A4(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n456_), .B(new_n772_), .C1(new_n812_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n297_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n800_), .A2(new_n604_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n802_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n808_), .A2(new_n806_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n811_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n595_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n814_), .A2(new_n817_), .A3(new_n819_), .A4(new_n821_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(KEYINPUT59), .A3(new_n456_), .A4(new_n772_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n827_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n297_), .A2(G113gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT118), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n825_), .B1(new_n837_), .B2(new_n839_), .ZN(G1340gat));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(KEYINPUT60), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n269_), .B2(KEYINPUT60), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT119), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n823_), .A2(new_n842_), .A3(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT120), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n269_), .B1(new_n827_), .B2(new_n836_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n841_), .B2(new_n847_), .ZN(G1341gat));
  INV_X1    g647(.A(G127gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n824_), .A2(new_n849_), .A3(new_n636_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n595_), .B1(new_n827_), .B2(new_n836_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n824_), .A2(new_n853_), .A3(new_n605_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n645_), .B1(new_n827_), .B2(new_n836_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n853_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT121), .B(new_n854_), .C1(new_n855_), .C2(new_n853_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1343gat));
  NOR4_X1   g659(.A1(new_n614_), .A2(new_n599_), .A3(new_n623_), .A4(new_n456_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n835_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n296_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n369_), .ZN(G1344gat));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n269_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n370_), .ZN(G1345gat));
  XNOR2_X1  g665(.A(KEYINPUT61), .B(G155gat), .ZN(new_n867_));
  INV_X1    g666(.A(new_n862_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n636_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT122), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n869_), .A2(KEYINPUT122), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n867_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n869_), .A2(KEYINPUT122), .ZN(new_n874_));
  INV_X1    g673(.A(new_n867_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n870_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(G1346gat));
  AOI21_X1  g676(.A(G162gat), .B1(new_n868_), .B2(new_n605_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n879_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n868_), .A2(G162gat), .A3(new_n580_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(G1347gat));
  NAND2_X1  g682(.A1(new_n614_), .A2(new_n403_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n632_), .A2(new_n884_), .A3(new_n296_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n318_), .B1(new_n835_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n886_), .A2(new_n887_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n812_), .A2(new_n822_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n525_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n626_), .A2(new_n403_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n297_), .A2(new_n460_), .ZN(new_n895_));
  OAI22_X1  g694(.A1(new_n889_), .A2(new_n890_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  OAI221_X1 g697(.A(KEYINPUT124), .B1(new_n894_), .B2(new_n895_), .C1(new_n889_), .C2(new_n890_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1348gat));
  INV_X1    g699(.A(new_n894_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n268_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n891_), .A2(new_n690_), .A3(new_n884_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n268_), .A2(G176gat), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n902_), .A2(new_n317_), .B1(new_n903_), .B2(new_n904_), .ZN(G1349gat));
  AOI21_X1  g704(.A(G183gat), .B1(new_n903_), .B2(new_n636_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n595_), .A2(new_n326_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n901_), .B2(new_n907_), .ZN(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n894_), .B2(new_n645_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n605_), .A2(new_n327_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n894_), .B2(new_n910_), .ZN(G1351gat));
  NAND2_X1  g710(.A1(new_n835_), .A2(new_n614_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n358_), .A2(new_n530_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n912_), .A2(new_n296_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  AOI21_X1  g714(.A(G197gat), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(KEYINPUT126), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918_));
  INV_X1    g717(.A(new_n913_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n892_), .A2(new_n297_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n920_), .B2(KEYINPUT125), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n916_), .B1(new_n917_), .B2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n405_), .B1(new_n920_), .B2(KEYINPUT125), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT126), .B1(new_n914_), .B2(new_n915_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n920_), .A2(KEYINPUT125), .A3(new_n918_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n922_), .A2(new_n926_), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n912_), .A2(new_n913_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n268_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g729(.A(KEYINPUT63), .B(G211gat), .Z(new_n931_));
  NAND3_X1  g730(.A1(new_n928_), .A2(new_n636_), .A3(new_n931_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n932_), .A2(KEYINPUT127), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(KEYINPUT127), .ZN(new_n934_));
  AOI211_X1 g733(.A(KEYINPUT63), .B(G211gat), .C1(new_n928_), .C2(new_n636_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(G1354gat));
  NAND3_X1  g735(.A1(new_n928_), .A2(new_n417_), .A3(new_n605_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n912_), .A2(new_n645_), .A3(new_n913_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n417_), .B2(new_n938_), .ZN(G1355gat));
endmodule


