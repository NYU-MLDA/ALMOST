//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_;
  XNOR2_X1  g000(.A(KEYINPUT74), .B(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G155gat), .B(G162gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(G141gat), .ZN(new_n207_));
  INV_X1    g006(.A(G148gat), .ZN(new_n208_));
  AOI22_X1  g007(.A1(new_n206_), .A2(KEYINPUT1), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n205_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n207_), .B(new_n208_), .C1(KEYINPUT83), .C2(KEYINPUT3), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n213_), .A2(new_n214_), .B1(KEYINPUT83), .B2(KEYINPUT3), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n205_), .B(KEYINPUT2), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n203_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n211_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G127gat), .B(G134gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(G113gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(G113gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n220_), .A2(G120gat), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(G120gat), .B1(new_n220_), .B2(new_n221_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  OAI22_X1  g024(.A1(new_n211_), .A2(new_n217_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT4), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT90), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G225gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT91), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT92), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n225_), .A2(new_n232_), .A3(KEYINPUT4), .A4(new_n226_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n226_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n228_), .A2(new_n231_), .A3(new_n233_), .A4(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n225_), .A2(new_n226_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n230_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT0), .B(G57gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G85gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(G1gat), .B(G29gat), .Z(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n237_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT98), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G8gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G15gat), .B(G22gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(G1gat), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT75), .ZN(new_n260_));
  INV_X1    g059(.A(G1gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n255_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n251_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(G8gat), .A3(new_n262_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT69), .B(G43gat), .ZN(new_n266_));
  INV_X1    g065(.A(G50gat), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n267_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G29gat), .B(G36gat), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n268_), .A2(new_n271_), .A3(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n273_), .A3(KEYINPUT78), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n264_), .A2(new_n265_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n250_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n264_), .A2(new_n265_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT15), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n268_), .A2(new_n271_), .A3(new_n269_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n271_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n273_), .A2(KEYINPUT15), .A3(new_n274_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n249_), .A3(new_n280_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n283_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G113gat), .B(G141gat), .ZN(new_n294_));
  INV_X1    g093(.A(G169gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(G197gat), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n283_), .A2(new_n292_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT8), .ZN(new_n303_));
  XOR2_X1   g102(.A(G85gat), .B(G92gat), .Z(new_n304_));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n305_));
  OAI22_X1  g104(.A1(new_n305_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(KEYINPUT7), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n305_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G99gat), .A2(G106gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n303_), .B(new_n304_), .C1(new_n308_), .C2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n306_), .A2(new_n307_), .ZN(new_n317_));
  AND3_X1   g116(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n320_), .A3(new_n309_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n303_), .B1(new_n321_), .B2(new_n304_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT67), .B1(new_n316_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G106gat), .ZN(new_n324_));
  INV_X1    g123(.A(G99gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT10), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT10), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G99gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT64), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT64), .B1(new_n326_), .B2(new_n328_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n324_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT65), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n304_), .A2(new_n332_), .A3(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n333_), .A2(new_n334_), .A3(G85gat), .A4(G92gat), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n331_), .A2(new_n336_), .A3(new_n337_), .A4(new_n320_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n304_), .B1(new_n308_), .B2(new_n314_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT8), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n315_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n323_), .A2(new_n338_), .A3(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G57gat), .B(G64gat), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT11), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(KEYINPUT11), .ZN(new_n346_));
  XOR2_X1   g145(.A(G71gat), .B(G78gat), .Z(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n346_), .A2(new_n347_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT12), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n343_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n338_), .B1(new_n316_), .B2(new_n322_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n350_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n351_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G230gat), .A2(G233gat), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n350_), .B(new_n338_), .C1(new_n322_), .C2(new_n316_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n353_), .A2(new_n357_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n359_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n358_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G120gat), .B(G148gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G204gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT5), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G176gat), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n364_), .A2(new_n368_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT13), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT68), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n371_), .B(KEYINPUT13), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT68), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(KEYINPUT23), .B2(new_n381_), .ZN(new_n383_));
  INV_X1    g182(.A(G176gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n295_), .A2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(KEYINPUT24), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT26), .B(G190gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n391_));
  AND2_X1   g190(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n385_), .A2(KEYINPUT24), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n383_), .A2(KEYINPUT80), .A3(new_n386_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT22), .B(G169gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n384_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n380_), .A2(new_n381_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n381_), .A2(KEYINPUT23), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n401_), .B(new_n394_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n399_), .A2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G71gat), .B(G99gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT30), .B(KEYINPUT31), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G15gat), .B(G43gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n224_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n413_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT94), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT27), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G211gat), .B(G218gat), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT21), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(KEYINPUT21), .ZN(new_n424_));
  XOR2_X1   g223(.A(G197gat), .B(G204gat), .Z(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n424_), .A2(new_n425_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n407_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n397_), .A2(KEYINPUT85), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n386_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT86), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n396_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n435_), .B(new_n386_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n430_), .A2(new_n432_), .A3(new_n434_), .A4(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n383_), .B1(G183gat), .B2(G190gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n400_), .B(KEYINPUT87), .Z(new_n439_));
  OAI211_X1 g238(.A(new_n438_), .B(new_n394_), .C1(G176gat), .C2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n428_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n429_), .A2(KEYINPUT20), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT19), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n437_), .A2(new_n440_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(new_n428_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n445_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n399_), .A2(new_n406_), .A3(new_n441_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G8gat), .B(G36gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n421_), .B1(new_n453_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n449_), .A2(new_n451_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n445_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n447_), .B1(new_n407_), .B2(new_n428_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n450_), .A3(new_n442_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n420_), .B1(new_n460_), .B2(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n450_), .B1(new_n463_), .B2(new_n442_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n459_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  AND4_X1   g268(.A1(new_n420_), .A2(new_n469_), .A3(new_n465_), .A4(KEYINPUT27), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT95), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n462_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n458_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n421_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G22gat), .B(G50gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT28), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n217_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n210_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n480_), .B2(KEYINPUT29), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n218_), .A2(new_n482_), .A3(new_n477_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT84), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(KEYINPUT29), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(new_n324_), .A3(new_n428_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490_));
  INV_X1    g289(.A(G78gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n324_), .B1(new_n487_), .B2(new_n428_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n492_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n487_), .A2(new_n428_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G106gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n497_), .B2(new_n488_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n486_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n492_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n486_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n484_), .A2(new_n485_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n495_), .A3(new_n488_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n505_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n471_), .A2(new_n472_), .A3(new_n475_), .A4(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n469_), .A2(new_n465_), .A3(KEYINPUT27), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT94), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n460_), .A2(new_n420_), .A3(new_n465_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n506_), .A2(new_n509_), .A3(new_n510_), .A4(new_n475_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT95), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n505_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT33), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n245_), .B(new_n515_), .ZN(new_n516_));
  OR3_X1    g315(.A1(new_n473_), .A2(new_n474_), .A3(KEYINPUT89), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT89), .B1(new_n473_), .B2(new_n474_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n228_), .A2(new_n230_), .A3(new_n233_), .A4(new_n236_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n519_), .A2(KEYINPUT93), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n238_), .A2(new_n231_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(KEYINPUT93), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n520_), .A2(new_n243_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .A4(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n458_), .A2(KEYINPUT32), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n453_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n462_), .A2(new_n464_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n247_), .B(new_n526_), .C1(new_n527_), .C2(new_n525_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n514_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n419_), .B1(new_n513_), .B2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n509_), .A2(new_n510_), .A3(new_n505_), .A4(new_n475_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT96), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n532_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n247_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n533_), .A2(new_n418_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  AOI211_X1 g335(.A(new_n302_), .B(new_n379_), .C1(new_n530_), .C2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G127gat), .B(G155gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G183gat), .B(G211gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n350_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n265_), .A3(new_n264_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n284_), .A2(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n542_), .B1(new_n548_), .B2(KEYINPUT17), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n542_), .A2(KEYINPUT17), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n548_), .A2(KEYINPUT77), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n343_), .A2(new_n290_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n354_), .A2(new_n275_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n557_), .A2(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT70), .B(G190gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(G218gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(G134gat), .B(G162gat), .Z(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(KEYINPUT36), .ZN(new_n568_));
  INV_X1    g367(.A(new_n562_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n554_), .A2(new_n569_), .A3(new_n560_), .A4(new_n559_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT71), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n563_), .A2(new_n573_), .A3(new_n568_), .A4(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n563_), .A2(new_n570_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n568_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n567_), .A2(KEYINPUT36), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(new_n576_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n568_), .B1(new_n563_), .B2(new_n570_), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n572_), .A2(new_n574_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(KEYINPUT73), .A3(new_n576_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n580_), .A2(KEYINPUT72), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT72), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n589_), .A3(new_n579_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n575_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT37), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n553_), .B1(new_n587_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n537_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT97), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n537_), .B2(new_n593_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n202_), .B(new_n248_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT38), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n553_), .A2(new_n585_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n537_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n535_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(G1324gat));
  INV_X1    g402(.A(KEYINPUT40), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n509_), .A2(new_n510_), .A3(new_n475_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n537_), .A2(new_n600_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(KEYINPUT99), .A2(KEYINPUT39), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(G8gat), .A3(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(KEYINPUT99), .A2(KEYINPUT39), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n610_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n607_), .A2(G8gat), .A3(new_n612_), .A4(new_n608_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n251_), .B(new_n606_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n605_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  AND4_X1   g415(.A1(new_n605_), .A2(new_n615_), .A3(new_n611_), .A4(new_n613_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n604_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n605_), .A3(new_n615_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n615_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n611_), .A2(new_n613_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT100), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n619_), .A2(new_n622_), .A3(KEYINPUT40), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n623_), .ZN(G1325gat));
  OAI21_X1  g423(.A(G15gat), .B1(new_n601_), .B2(new_n419_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT41), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n594_), .A2(G15gat), .A3(new_n419_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(G1326gat));
  OAI21_X1  g427(.A(G22gat), .B1(new_n601_), .B2(new_n505_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT101), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n631_), .ZN(new_n633_));
  OR3_X1    g432(.A1(new_n594_), .A2(G22gat), .A3(new_n505_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(G1327gat));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n530_), .A2(new_n536_), .ZN(new_n637_));
  AND4_X1   g436(.A1(KEYINPUT73), .A2(new_n575_), .A3(new_n576_), .A4(new_n580_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT73), .B1(new_n585_), .B2(new_n576_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n592_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n637_), .B2(new_n641_), .ZN(new_n642_));
  AOI211_X1 g441(.A(KEYINPUT43), .B(new_n640_), .C1(new_n530_), .C2(new_n536_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n553_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n379_), .A2(new_n645_), .A3(new_n302_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n642_), .A2(new_n643_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n646_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n647_), .A2(new_n248_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n653_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(G29gat), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n585_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n530_), .B2(new_n536_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n646_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n535_), .A2(G29gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(G1328gat));
  NAND2_X1  g460(.A1(new_n647_), .A2(new_n651_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n606_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G36gat), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  OR3_X1    g463(.A1(new_n659_), .A2(G36gat), .A3(new_n663_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT45), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(KEYINPUT45), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n664_), .B(KEYINPUT46), .C1(new_n667_), .C2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1329gat));
  INV_X1    g472(.A(KEYINPUT47), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n647_), .A2(new_n651_), .A3(G43gat), .A4(new_n418_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  INV_X1    g475(.A(G43gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n659_), .B2(new_n419_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n676_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n676_), .B1(new_n675_), .B2(new_n678_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n674_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n681_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(KEYINPUT47), .A3(new_n679_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1330gat));
  OAI21_X1  g484(.A(G50gat), .B1(new_n662_), .B2(new_n505_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n514_), .A2(new_n267_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT104), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n659_), .B2(new_n688_), .ZN(G1331gat));
  AOI211_X1 g488(.A(new_n301_), .B(new_n378_), .C1(new_n530_), .C2(new_n536_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n593_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G57gat), .B1(new_n692_), .B2(new_n248_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n600_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n535_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(G57gat), .B2(new_n695_), .ZN(G1332gat));
  OAI21_X1  g495(.A(G64gat), .B1(new_n694_), .B2(new_n663_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT48), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n691_), .A2(G64gat), .A3(new_n663_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT105), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n694_), .B2(new_n419_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n419_), .A2(G71gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n691_), .B2(new_n704_), .ZN(G1334gat));
  OAI21_X1  g504(.A(G78gat), .B1(new_n694_), .B2(new_n505_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT50), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n706_), .B(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n692_), .A2(new_n491_), .A3(new_n514_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1335gat));
  NOR3_X1   g510(.A1(new_n378_), .A2(new_n645_), .A3(new_n301_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n658_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n248_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n644_), .A2(new_n712_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n247_), .A2(G85gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT108), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n714_), .B1(new_n715_), .B2(new_n717_), .ZN(G1336gat));
  AOI21_X1  g517(.A(G92gat), .B1(new_n713_), .B2(new_n606_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n606_), .A2(G92gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n715_), .B2(new_n720_), .ZN(G1337gat));
  NAND2_X1  g520(.A1(new_n715_), .A2(new_n418_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G99gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n713_), .B(new_n418_), .C1(new_n330_), .C2(new_n329_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n724_), .A3(new_n727_), .ZN(new_n728_));
  OR2_X1    g527(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(G1338gat));
  OAI211_X1 g529(.A(new_n514_), .B(new_n712_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G106gat), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n713_), .A2(KEYINPUT111), .A3(new_n324_), .A4(new_n514_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n658_), .A2(new_n324_), .A3(new_n712_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(new_n505_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n735_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT112), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n734_), .A2(new_n743_), .A3(new_n735_), .A4(new_n740_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n742_), .A2(KEYINPUT53), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT53), .B1(new_n742_), .B2(new_n744_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1339gat));
  NAND4_X1  g546(.A1(new_n533_), .A2(new_n418_), .A3(new_n534_), .A4(new_n248_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n371_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n249_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n291_), .A2(new_n250_), .A3(new_n280_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n297_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n300_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n750_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n370_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n360_), .A2(KEYINPUT115), .ZN(new_n758_));
  INV_X1    g557(.A(new_n359_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n358_), .A4(new_n353_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n760_), .A2(new_n353_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n362_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n358_), .B1(new_n760_), .B2(new_n353_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n758_), .B(new_n762_), .C1(new_n768_), .C2(new_n764_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n769_), .A4(new_n368_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n301_), .B(new_n757_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n767_), .A2(new_n368_), .A3(new_n769_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n771_), .A3(new_n770_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n756_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT117), .B1(new_n778_), .B2(new_n585_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n776_), .A2(new_n771_), .A3(new_n770_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n755_), .B1(new_n780_), .B2(new_n772_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n657_), .ZN(new_n783_));
  XOR2_X1   g582(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n776_), .A2(new_n770_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n757_), .A3(new_n754_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n641_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n781_), .A2(KEYINPUT57), .A3(new_n657_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n781_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n657_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n785_), .A2(new_n789_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n794_), .A2(new_n553_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n376_), .A2(new_n301_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n640_), .A2(new_n645_), .A3(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(KEYINPUT113), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(KEYINPUT113), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AOI211_X1 g602(.A(KEYINPUT114), .B(KEYINPUT54), .C1(new_n797_), .C2(KEYINPUT113), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n593_), .B2(new_n796_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT114), .B1(new_n807_), .B2(KEYINPUT54), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n801_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n798_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n805_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n749_), .B1(new_n795_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n794_), .A2(new_n553_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(new_n810_), .A3(new_n805_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(KEYINPUT59), .A3(new_n749_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(G113gat), .B(new_n301_), .C1(new_n815_), .C2(new_n819_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n817_), .A2(KEYINPUT120), .A3(new_n749_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT120), .B1(new_n817_), .B2(new_n749_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n302_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n820_), .B1(new_n825_), .B2(G113gat), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(G1340gat));
  INV_X1    g626(.A(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n378_), .B2(KEYINPUT60), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n828_), .A2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n829_), .B(new_n830_), .C1(new_n821_), .C2(new_n823_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n378_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n828_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT121), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n831_), .B(new_n835_), .C1(new_n832_), .C2(new_n828_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1341gat));
  OAI211_X1 g636(.A(G127gat), .B(new_n645_), .C1(new_n815_), .C2(new_n819_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n553_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(G127gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n842_), .B(new_n585_), .C1(new_n821_), .C2(new_n823_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n640_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT122), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n843_), .B(new_n847_), .C1(new_n844_), .C2(new_n842_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1343gat));
  NAND4_X1  g648(.A1(new_n419_), .A2(new_n514_), .A3(new_n663_), .A4(new_n248_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT123), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n817_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n302_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n207_), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n378_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n208_), .ZN(G1345gat));
  NOR2_X1   g655(.A1(new_n852_), .A2(new_n553_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT61), .B(G155gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  INV_X1    g658(.A(new_n852_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n860_), .A2(G162gat), .A3(new_n641_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G162gat), .B1(new_n860_), .B2(new_n585_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n862_), .A2(KEYINPUT124), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(KEYINPUT124), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n863_), .B2(new_n864_), .ZN(G1347gat));
  NOR3_X1   g664(.A1(new_n419_), .A2(new_n663_), .A3(new_n248_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n817_), .A2(new_n505_), .A3(new_n301_), .A4(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G169gat), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n867_), .A2(new_n439_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n870_), .A2(new_n871_), .A3(KEYINPUT125), .A4(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1348gat));
  NOR2_X1   g676(.A1(KEYINPUT126), .A2(G176gat), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n817_), .A2(new_n505_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n379_), .A3(new_n866_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(KEYINPUT126), .A2(G176gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n880_), .B2(new_n878_), .ZN(G1349gat));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n866_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI211_X1 g684(.A(KEYINPUT127), .B(G183gat), .C1(new_n885_), .C2(new_n645_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(KEYINPUT127), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n884_), .A2(new_n553_), .A3(new_n392_), .A4(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1350gat));
  OAI21_X1  g688(.A(G190gat), .B1(new_n884_), .B2(new_n640_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n585_), .A2(new_n390_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n884_), .B2(new_n891_), .ZN(G1351gat));
  NAND2_X1  g691(.A1(new_n817_), .A2(new_n535_), .ZN(new_n893_));
  NOR4_X1   g692(.A1(new_n893_), .A2(new_n418_), .A3(new_n505_), .A4(new_n663_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n301_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n379_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n645_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT63), .B(G211gat), .Z(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n899_), .B2(new_n901_), .ZN(G1354gat));
  AOI21_X1  g701(.A(G218gat), .B1(new_n894_), .B2(new_n585_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n894_), .A2(G218gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n641_), .B2(new_n904_), .ZN(G1355gat));
endmodule


