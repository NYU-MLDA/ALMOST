//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G127gat), .ZN(new_n204_));
  INV_X1    g003(.A(G127gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G134gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT85), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT85), .B1(new_n204_), .B2(new_n206_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n206_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT85), .ZN(new_n213_));
  INV_X1    g012(.A(new_n202_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n209_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222_));
  AND3_X1   g021(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT87), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT1), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n221_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n217_), .B(KEYINPUT2), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n219_), .A2(KEYINPUT88), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n219_), .A2(KEYINPUT88), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT3), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n233_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n216_), .A2(new_n235_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n209_), .A2(new_n215_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT88), .ZN(new_n247_));
  NOR4_X1   g046(.A1(new_n247_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n237_), .B1(new_n219_), .B2(KEYINPUT88), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n242_), .B1(new_n250_), .B2(new_n236_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n246_), .B1(new_n234_), .B2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G225gat), .A2(G233gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n246_), .B(new_n256_), .C1(new_n234_), .C2(new_n251_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n254_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n245_), .A2(KEYINPUT4), .A3(new_n252_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT96), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n255_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT0), .ZN(new_n266_));
  INV_X1    g065(.A(G57gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(G85gat), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n271_), .B(new_n255_), .C1(new_n263_), .C2(new_n262_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT18), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G204gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G197gat), .ZN(new_n280_));
  INV_X1    g079(.A(G197gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G204gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT21), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(KEYINPUT90), .A3(new_n283_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n281_), .B2(G204gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n282_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n280_), .A2(new_n290_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT21), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT91), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT91), .ZN(new_n297_));
  INV_X1    g096(.A(G211gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(G218gat), .ZN(new_n299_));
  INV_X1    g098(.A(G218gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(G211gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n297_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n289_), .A2(new_n294_), .A3(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n296_), .A2(new_n302_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n287_), .A2(new_n283_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n310_), .A2(KEYINPUT80), .A3(G183gat), .A4(G190gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(G183gat), .A3(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT80), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(KEYINPUT23), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n311_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n319_), .A2(KEYINPUT24), .ZN(new_n320_));
  INV_X1    g119(.A(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n318_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n325_));
  INV_X1    g124(.A(G183gat), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n325_), .A2(new_n326_), .A3(KEYINPUT25), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT25), .B(G183gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G190gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT79), .B1(new_n330_), .B2(KEYINPUT26), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G190gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(KEYINPUT79), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n317_), .B(new_n324_), .C1(new_n329_), .C2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n321_), .B2(KEYINPUT22), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT81), .B(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n321_), .A2(KEYINPUT81), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n321_), .A2(KEYINPUT81), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n335_), .B(KEYINPUT22), .C1(new_n340_), .C2(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n339_), .A2(new_n322_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n315_), .A2(KEYINPUT23), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n312_), .A3(KEYINPUT83), .ZN(new_n345_));
  OR3_X1    g144(.A1(new_n315_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n326_), .A2(new_n330_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n319_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n334_), .B1(new_n343_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT84), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n339_), .A2(new_n322_), .A3(new_n342_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n348_), .A3(new_n319_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT84), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n334_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n309_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n317_), .A2(new_n347_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G169gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT94), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n319_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(KEYINPUT94), .A2(G169gat), .A3(G176gat), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n361_), .A2(new_n322_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n328_), .A2(new_n332_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n324_), .A2(new_n367_), .A3(new_n346_), .A4(new_n345_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT20), .B1(new_n308_), .B2(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n356_), .A2(new_n359_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n359_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n351_), .A2(new_n355_), .A3(new_n309_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT20), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n308_), .B2(new_n369_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n278_), .B1(new_n371_), .B2(new_n376_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n371_), .A2(new_n376_), .A3(new_n278_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(KEYINPUT95), .ZN(new_n379_));
  INV_X1    g178(.A(new_n278_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n373_), .A2(new_n375_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n359_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n355_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n354_), .B1(new_n353_), .B2(new_n334_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n308_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n370_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n372_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n380_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT27), .B1(new_n379_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n382_), .A2(new_n380_), .A3(new_n387_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT27), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT97), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n351_), .A2(new_n355_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n370_), .B1(new_n395_), .B2(new_n308_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n396_), .B2(new_n372_), .ZN(new_n397_));
  OAI211_X1 g196(.A(KEYINPUT97), .B(new_n359_), .C1(new_n356_), .C2(new_n370_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n397_), .B(new_n398_), .C1(new_n359_), .C2(new_n381_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n393_), .B1(new_n399_), .B2(new_n278_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n391_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n395_), .A2(KEYINPUT30), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G71gat), .B(G99gat), .ZN(new_n404_));
  INV_X1    g203(.A(G43gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407_));
  INV_X1    g206(.A(G15gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n406_), .B(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n395_), .A2(KEYINPUT30), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n403_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n403_), .B2(new_n411_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n402_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n216_), .B(KEYINPUT31), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n414_), .B(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n232_), .B1(new_n225_), .B2(new_n230_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n244_), .B1(new_n418_), .B2(new_n221_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(KEYINPUT29), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT28), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT29), .B1(new_n234_), .B2(new_n251_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT92), .B1(G228gat), .B2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(KEYINPUT92), .A2(G228gat), .A3(G233gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n424_), .A2(new_n308_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n424_), .B2(new_n308_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n423_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n424_), .A2(new_n308_), .A3(new_n428_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n419_), .A2(KEYINPUT29), .B1(new_n304_), .B2(new_n307_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n432_), .B(new_n422_), .C1(new_n433_), .C2(new_n426_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G22gat), .B(G50gat), .Z(new_n435_));
  AND3_X1   g234(.A1(new_n431_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n421_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n435_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n429_), .A2(new_n430_), .A3(new_n423_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n424_), .A2(new_n308_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n425_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n422_), .B1(new_n442_), .B2(new_n432_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n439_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n421_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n431_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  AND4_X1   g247(.A1(new_n274_), .A2(new_n401_), .A3(new_n417_), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT27), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n388_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n377_), .A2(KEYINPUT95), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n438_), .A2(new_n447_), .A3(new_n270_), .A4(new_n272_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n398_), .B1(new_n359_), .B2(new_n381_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n385_), .A2(new_n386_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT97), .B1(new_n457_), .B2(new_n359_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(KEYINPUT27), .B(new_n392_), .C1(new_n459_), .C2(new_n380_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n453_), .A2(new_n455_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT98), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT98), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n453_), .A2(new_n455_), .A3(new_n463_), .A4(new_n460_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n382_), .A2(new_n387_), .A3(new_n465_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n273_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n379_), .A2(new_n390_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n272_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n263_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(KEYINPUT33), .A3(new_n255_), .A4(new_n271_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n260_), .A2(new_n254_), .A3(new_n257_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n253_), .A2(new_n258_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n269_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n472_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n469_), .B1(new_n470_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n448_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n462_), .A2(new_n464_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n417_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n449_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT72), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G120gat), .B(G148gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT5), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT71), .ZN(new_n489_));
  XOR2_X1   g288(.A(G176gat), .B(G204gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G71gat), .B(G78gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(KEYINPUT11), .B2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT68), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n495_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n497_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT69), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G99gat), .ZN(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n507_), .B(new_n508_), .C1(new_n509_), .C2(KEYINPUT67), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n510_), .B1(new_n511_), .B2(KEYINPUT7), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n509_), .A2(new_n507_), .A3(new_n508_), .A4(KEYINPUT67), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G85gat), .B(G92gat), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(KEYINPUT8), .A3(new_n515_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(KEYINPUT65), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n520_), .A2(new_n521_), .A3(KEYINPUT65), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT64), .B(G85gat), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n522_), .B(new_n523_), .C1(new_n526_), .C2(KEYINPUT9), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT10), .B(G99gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n508_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n506_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n518_), .A2(new_n519_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n500_), .A2(new_n501_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n496_), .A2(new_n497_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n503_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT12), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G230gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n531_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n535_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n534_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n532_), .A2(new_n533_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(new_n537_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n531_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n538_), .A2(new_n539_), .A3(new_n543_), .A4(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n503_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n531_), .B1(new_n503_), .B2(new_n535_), .ZN(new_n549_));
  OAI211_X1 g348(.A(G230gat), .B(G233gat), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT70), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n486_), .B(new_n492_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n491_), .B1(new_n556_), .B2(new_n552_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n547_), .A2(new_n550_), .A3(new_n491_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT72), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n555_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n562_), .A2(KEYINPUT13), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(KEYINPUT13), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n492_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(KEYINPUT72), .B2(new_n559_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n567_), .A2(new_n562_), .A3(KEYINPUT13), .A4(new_n555_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G29gat), .B(G36gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(G43gat), .B(G50gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n572_), .B(KEYINPUT15), .Z(new_n573_));
  INV_X1    g372(.A(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(G8gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(G22gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(G15gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n408_), .A2(G22gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT75), .ZN(new_n581_));
  XOR2_X1   g380(.A(G1gat), .B(G8gat), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n580_), .A2(KEYINPUT75), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(KEYINPUT75), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n582_), .A3(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n573_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n587_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n572_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n572_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n596_), .A2(G229gat), .A3(G233gat), .A4(new_n592_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n595_), .A2(new_n597_), .A3(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT77), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n485_), .A2(new_n569_), .A3(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n609_));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT35), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n531_), .B2(new_n572_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n531_), .B2(new_n573_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n611_), .A2(new_n612_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(KEYINPUT36), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n620_), .B(KEYINPUT36), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n617_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT37), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n590_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(new_n544_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G127gat), .B(G155gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n534_), .B1(new_n634_), .B2(KEYINPUT17), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n629_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n629_), .A2(new_n635_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n634_), .A2(KEYINPUT17), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n626_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n608_), .A2(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n641_), .A2(G1gat), .A3(new_n274_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n643_));
  XOR2_X1   g442(.A(new_n642_), .B(new_n643_), .Z(new_n644_));
  INV_X1    g443(.A(new_n605_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n569_), .A2(new_n645_), .A3(new_n639_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n485_), .A2(new_n625_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT100), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n574_), .B1(new_n649_), .B2(new_n273_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n644_), .A2(new_n650_), .ZN(G1324gat));
  INV_X1    g450(.A(new_n641_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n401_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n575_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n646_), .A2(new_n647_), .A3(new_n653_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G8gat), .B1(new_n655_), .B2(new_n656_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT39), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT39), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n654_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT40), .B(new_n654_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  AOI21_X1  g465(.A(new_n408_), .B1(new_n649_), .B2(new_n417_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n652_), .A2(new_n408_), .A3(new_n417_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(new_n448_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n577_), .B1(new_n649_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT42), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n652_), .A2(new_n577_), .A3(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1327gat));
  NAND4_X1  g476(.A1(new_n565_), .A2(new_n568_), .A3(new_n605_), .A4(new_n639_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n482_), .A2(new_n464_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n391_), .A2(new_n454_), .A3(new_n400_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n463_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n484_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n449_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n680_), .B1(new_n686_), .B2(new_n626_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT37), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n625_), .B(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n485_), .A2(KEYINPUT43), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n679_), .B1(new_n687_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n485_), .B2(new_n689_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n682_), .A2(new_n463_), .B1(new_n448_), .B2(new_n481_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n417_), .B1(new_n695_), .B2(new_n462_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n680_), .B(new_n626_), .C1(new_n696_), .C2(new_n449_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n678_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT44), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n693_), .A2(new_n273_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(G29gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n625_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n639_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n608_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n273_), .A2(new_n701_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT102), .ZN(new_n707_));
  OAI22_X1  g506(.A1(new_n700_), .A2(new_n701_), .B1(new_n705_), .B2(new_n707_), .ZN(G1328gat));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n653_), .B1(new_n698_), .B2(KEYINPUT44), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n692_), .B(new_n678_), .C1(new_n694_), .C2(new_n697_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G36gat), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n569_), .A2(new_n607_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n401_), .A2(G36gat), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n713_), .A2(new_n686_), .A3(new_n704_), .A4(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT45), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n712_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT46), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n709_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n719_), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT104), .B(new_n721_), .C1(new_n712_), .C2(new_n716_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n718_), .A2(KEYINPUT46), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n720_), .A2(new_n722_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n715_), .B(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n693_), .A2(new_n653_), .A3(new_n699_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(G36gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT104), .B1(new_n729_), .B2(new_n721_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n717_), .A2(new_n709_), .A3(new_n719_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n723_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n725_), .A2(new_n732_), .ZN(G1329gat));
  OAI21_X1  g532(.A(new_n405_), .B1(new_n705_), .B2(new_n484_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n693_), .A2(G43gat), .A3(new_n417_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n711_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g536(.A1(new_n693_), .A2(G50gat), .A3(new_n673_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n705_), .A2(new_n448_), .ZN(new_n739_));
  OAI22_X1  g538(.A1(new_n738_), .A2(new_n711_), .B1(G50gat), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT105), .Z(G1331gat));
  NOR2_X1   g540(.A1(new_n606_), .A2(new_n639_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n647_), .A2(new_n569_), .A3(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT106), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n274_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n569_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n485_), .A3(new_n605_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n640_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n746_), .A2(new_n751_), .ZN(G1332gat));
  INV_X1    g551(.A(G64gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n753_), .A3(new_n653_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n744_), .A2(new_n653_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G64gat), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT48), .B(new_n753_), .C1(new_n744_), .C2(new_n653_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(KEYINPUT107), .B(new_n754_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1333gat));
  OR3_X1    g562(.A1(new_n749_), .A2(G71gat), .A3(new_n484_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G71gat), .B1(new_n745_), .B2(new_n484_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(KEYINPUT49), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(KEYINPUT49), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n764_), .B1(new_n766_), .B2(new_n767_), .ZN(G1334gat));
  OAI21_X1  g567(.A(G78gat), .B1(new_n745_), .B2(new_n448_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT50), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n448_), .A2(G78gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n749_), .B2(new_n771_), .ZN(G1335gat));
  AND2_X1   g571(.A1(new_n748_), .A2(new_n704_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n273_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n569_), .A2(new_n645_), .A3(new_n639_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT108), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n274_), .A2(new_n524_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n525_), .A3(new_n653_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n777_), .A2(new_n653_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n525_), .ZN(G1337gat));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n528_), .A3(new_n417_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n776_), .A2(new_n417_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n507_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n785_), .B(new_n786_), .Z(G1338gat));
  NAND3_X1  g586(.A1(new_n773_), .A2(new_n508_), .A3(new_n673_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n776_), .A2(new_n673_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n508_), .B1(new_n790_), .B2(KEYINPUT110), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n791_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n788_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n788_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  NAND2_X1  g600(.A1(new_n417_), .A2(new_n448_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n653_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n538_), .A2(KEYINPUT55), .A3(new_n543_), .A4(new_n546_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(G230gat), .A4(G233gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n549_), .B1(new_n531_), .B2(new_n545_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(G230gat), .A3(G233gat), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(KEYINPUT55), .A3(new_n538_), .A4(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n547_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n808_), .A2(new_n811_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n492_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n492_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n558_), .A2(new_n605_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT112), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n596_), .A2(new_n592_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n602_), .B1(new_n822_), .B2(new_n594_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n593_), .A2(new_n594_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n825_), .A2(new_n827_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n819_), .A2(new_n821_), .B1(new_n561_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n805_), .B1(new_n829_), .B2(new_n625_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n828_), .A2(new_n831_), .A3(new_n558_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n828_), .B2(new_n558_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n818_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT56), .B1(new_n814_), .B2(new_n492_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n834_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n626_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n820_), .B(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n828_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n567_), .B2(new_n555_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT57), .B(new_n702_), .C1(new_n844_), .C2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n830_), .A2(new_n841_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n639_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n850_));
  NAND4_X1  g649(.A1(new_n747_), .A2(new_n689_), .A3(new_n742_), .A4(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n850_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n689_), .A2(new_n742_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n569_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n274_), .B(new_n804_), .C1(new_n849_), .C2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(G113gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n605_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(KEYINPUT116), .A3(KEYINPUT59), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n849_), .A2(new_n855_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(KEYINPUT116), .A3(new_n273_), .A4(new_n803_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n607_), .B1(new_n859_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n858_), .B1(new_n864_), .B2(new_n857_), .ZN(G1340gat));
  XNOR2_X1  g664(.A(KEYINPUT117), .B(G120gat), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n747_), .A2(KEYINPUT60), .A3(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n867_), .A2(KEYINPUT60), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n856_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT59), .B1(new_n856_), .B2(KEYINPUT116), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n861_), .A2(new_n862_), .ZN(new_n872_));
  OAI211_X1 g671(.A(KEYINPUT118), .B(new_n569_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n867_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n859_), .A2(new_n863_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT118), .B1(new_n875_), .B2(new_n569_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n870_), .B1(new_n874_), .B2(new_n876_), .ZN(G1341gat));
  AOI21_X1  g676(.A(G127gat), .B1(new_n856_), .B2(new_n703_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT119), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n639_), .A2(new_n205_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n875_), .B2(new_n880_), .ZN(G1342gat));
  AOI21_X1  g680(.A(G134gat), .B1(new_n856_), .B2(new_n625_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT120), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT121), .B(G134gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n689_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n875_), .B2(new_n885_), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n860_), .A2(new_n273_), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n887_), .A2(new_n417_), .A3(new_n448_), .A4(new_n653_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n605_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT122), .B(G141gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n569_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n888_), .A2(new_n703_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n888_), .A2(new_n897_), .A3(new_n625_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n888_), .A2(new_n626_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1347gat));
  NOR3_X1   g699(.A1(new_n802_), .A2(new_n273_), .A3(new_n401_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n860_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n605_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(G169gat), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n903_), .B2(G169gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  AOI211_X1 g707(.A(KEYINPUT124), .B(new_n904_), .C1(new_n903_), .C2(G169gat), .ZN(new_n909_));
  INV_X1    g708(.A(new_n361_), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n908_), .A2(new_n909_), .B1(new_n910_), .B2(new_n903_), .ZN(G1348gat));
  NAND2_X1  g710(.A1(new_n902_), .A2(new_n569_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g712(.A1(new_n902_), .A2(new_n703_), .ZN(new_n914_));
  MUX2_X1   g713(.A(new_n328_), .B(G183gat), .S(new_n914_), .Z(G1350gat));
  NAND3_X1  g714(.A1(new_n902_), .A2(new_n625_), .A3(new_n332_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n902_), .A2(new_n626_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n330_), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n401_), .A2(new_n417_), .A3(new_n454_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n860_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT125), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n860_), .A2(new_n922_), .A3(new_n919_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n605_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n569_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  AND2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n924_), .B(new_n703_), .C1(new_n929_), .C2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n924_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n639_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n933_), .B2(new_n929_), .ZN(G1354gat));
  NOR3_X1   g733(.A1(new_n932_), .A2(new_n300_), .A3(new_n689_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n702_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  AOI21_X1  g736(.A(G218gat), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  OR2_X1    g737(.A1(new_n936_), .A2(new_n937_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n935_), .B1(new_n938_), .B2(new_n939_), .ZN(G1355gat));
endmodule


