//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n203_), .B1(new_n204_), .B2(new_n202_), .ZN(new_n205_));
  OR3_X1    g004(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n205_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT25), .ZN(new_n214_));
  OR2_X1    g013(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n213_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n222_));
  OAI211_X1 g021(.A(G183gat), .B(G190gat), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n202_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n215_), .A2(new_n216_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n223_), .B(new_n225_), .C1(G190gat), .C2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G169gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n220_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT30), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT31), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT83), .B(G15gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n241_), .A2(new_n242_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n243_), .B(new_n244_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT85), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G127gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(G134gat), .ZN(new_n250_));
  INV_X1    g049(.A(G134gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(G127gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT85), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G113gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(G120gat), .ZN(new_n256_));
  INV_X1    g055(.A(G120gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(G113gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT86), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(G113gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(G120gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT86), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n254_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n248_), .A2(new_n253_), .A3(new_n259_), .A4(new_n263_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT87), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268_));
  AND4_X1   g067(.A1(new_n248_), .A2(new_n253_), .A3(new_n259_), .A4(new_n263_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n248_), .A2(new_n253_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n245_), .A2(new_n267_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n245_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n267_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n236_), .A2(new_n272_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n272_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n235_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n280_));
  INV_X1    g079(.A(G197gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(G204gat), .A3(new_n283_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n281_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT91), .B1(new_n281_), .B2(G204gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G218gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G211gat), .ZN(new_n289_));
  INV_X1    g088(.A(G211gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G218gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n291_), .A3(KEYINPUT92), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT92), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n290_), .A2(G218gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n288_), .A2(G211gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n287_), .A2(KEYINPUT21), .A3(new_n292_), .A4(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT21), .ZN(new_n298_));
  INV_X1    g097(.A(G204gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(G197gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n299_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n303_), .B2(KEYINPUT90), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n305_), .B(new_n299_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n298_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n296_), .A2(new_n292_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n284_), .A2(new_n285_), .A3(new_n298_), .A4(new_n286_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n297_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n229_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT95), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n313_), .B1(new_n205_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n202_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n224_), .A2(G183gat), .A3(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n314_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT95), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n312_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n211_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT25), .B(G183gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n213_), .A2(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n322_), .A2(new_n223_), .A3(new_n225_), .A4(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n311_), .B1(new_n321_), .B2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(G204gat), .B1(new_n282_), .B2(new_n283_), .ZN(new_n328_));
  OAI22_X1  g127(.A1(new_n328_), .A2(new_n305_), .B1(G197gat), .B2(new_n299_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n306_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT21), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n308_), .A2(new_n309_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n212_), .A2(new_n219_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n297_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n327_), .A2(KEYINPUT20), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT98), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT95), .B1(new_n318_), .B2(new_n319_), .ZN(new_n341_));
  AOI211_X1 g140(.A(new_n313_), .B(new_n314_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n229_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n333_), .A2(new_n343_), .A3(new_n297_), .A4(new_n325_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n311_), .A2(new_n231_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n338_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n344_), .A2(KEYINPUT20), .A3(new_n345_), .A4(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n339_), .A2(new_n340_), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT20), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n343_), .A2(new_n325_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(new_n311_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n346_), .B1(new_n358_), .B2(new_n335_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n347_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n340_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n344_), .A2(KEYINPUT20), .A3(new_n345_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n338_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n346_), .A3(new_n335_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(KEYINPUT32), .A4(new_n353_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n355_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT2), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n369_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G155gat), .B(G162gat), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G155gat), .ZN(new_n378_));
  INV_X1    g177(.A(G162gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT1), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT1), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(G155gat), .A3(G162gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n379_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G141gat), .B(G148gat), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n377_), .A2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n266_), .B2(new_n265_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT88), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n377_), .A2(new_n386_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n377_), .B2(new_n386_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n274_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396_));
  AOI211_X1 g195(.A(new_n396_), .B(new_n388_), .C1(new_n274_), .C2(new_n392_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n267_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT87), .B1(new_n265_), .B2(new_n266_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n392_), .B(new_n396_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n394_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n395_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n395_), .B(new_n407_), .C1(new_n397_), .C2(new_n402_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(KEYINPUT99), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n403_), .A2(new_n412_), .A3(new_n408_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n366_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(KEYINPUT97), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT33), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n410_), .A2(KEYINPUT97), .A3(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n395_), .A2(new_n396_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n400_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n408_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n416_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n352_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n339_), .A2(new_n353_), .A3(new_n347_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT96), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n426_), .B(new_n352_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n414_), .B1(new_n422_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n392_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n432_), .B(new_n311_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n387_), .A2(KEYINPUT29), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT93), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT93), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n387_), .A2(new_n438_), .A3(KEYINPUT29), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n311_), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(G228gat), .A3(G233gat), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n431_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n441_), .A3(new_n431_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n392_), .A2(KEYINPUT29), .ZN(new_n446_));
  XOR2_X1   g245(.A(G22gat), .B(G50gat), .Z(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(KEYINPUT28), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n446_), .B(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n442_), .B2(KEYINPUT94), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n445_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n443_), .A2(KEYINPUT94), .A3(new_n444_), .A4(new_n449_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n429_), .A2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n451_), .A2(new_n452_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n424_), .A2(KEYINPUT27), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n352_), .B(KEYINPUT100), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT101), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n363_), .A2(new_n364_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n457_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT101), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT27), .A4(new_n424_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n411_), .A2(new_n413_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n425_), .A2(new_n467_), .A3(new_n427_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n455_), .A2(new_n465_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n279_), .B1(new_n454_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n279_), .A2(new_n466_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n465_), .A2(new_n453_), .A3(new_n468_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT102), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT102), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n465_), .A2(new_n453_), .A3(new_n474_), .A4(new_n468_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n471_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G113gat), .B(G141gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G169gat), .B(G197gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT74), .B(G1gat), .Z(new_n481_));
  INV_X1    g280(.A(G8gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT73), .B(G15gat), .ZN(new_n484_));
  INV_X1    g283(.A(G22gat), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n485_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G1gat), .B(G8gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n483_), .A2(new_n486_), .A3(new_n487_), .A4(new_n489_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G29gat), .B(G36gat), .Z(new_n494_));
  XOR2_X1   g293(.A(G43gat), .B(G50gat), .Z(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n493_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(KEYINPUT15), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n494_), .B(new_n495_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n499_), .A2(new_n502_), .A3(new_n492_), .A4(new_n491_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT78), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n493_), .A2(new_n500_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n498_), .ZN(new_n507_));
  OAI221_X1 g306(.A(new_n480_), .B1(new_n497_), .B2(new_n498_), .C1(new_n505_), .C2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n480_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n499_), .A2(new_n502_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n491_), .A2(new_n492_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n504_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n503_), .A2(KEYINPUT78), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n507_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n497_), .A2(new_n498_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n509_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n508_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT79), .B(new_n509_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT80), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n477_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G85gat), .B(G92gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n526_), .B2(KEYINPUT8), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT6), .Z(new_n529_));
  NOR2_X1   g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n527_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n526_), .A2(KEYINPUT8), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n527_), .B(new_n534_), .C1(new_n529_), .C2(new_n532_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT9), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n525_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT10), .B(G99gat), .Z(new_n541_));
  INV_X1    g340(.A(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(G85gat), .A3(G92gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n528_), .B(KEYINPUT6), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n540_), .A2(new_n543_), .A3(new_n544_), .A4(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n538_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  OAI22_X1  g348(.A1(new_n547_), .A2(new_n496_), .B1(KEYINPUT35), .B2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n547_), .B2(new_n510_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n551_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G190gat), .B(G218gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT70), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT71), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n554_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n557_), .B(KEYINPUT36), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n554_), .A2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n524_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n554_), .A2(new_n561_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n567_), .B(new_n523_), .C1(new_n554_), .C2(new_n564_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT64), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT66), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT11), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n573_), .A2(KEYINPUT66), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT11), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(KEYINPUT66), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n575_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n574_), .A2(KEYINPUT11), .A3(new_n580_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n546_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n572_), .B1(new_n587_), .B2(KEYINPUT67), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(KEYINPUT67), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n586_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n588_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n584_), .A2(KEYINPUT68), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT68), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n582_), .A2(new_n583_), .A3(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n595_), .A2(KEYINPUT12), .A3(new_n547_), .A4(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT69), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n590_), .B2(new_n572_), .ZN(new_n600_));
  AOI211_X1 g399(.A(KEYINPUT69), .B(new_n571_), .C1(new_n584_), .C2(new_n586_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n594_), .B(new_n598_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT5), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n592_), .A2(new_n602_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n592_), .B2(new_n602_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT13), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT13), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n511_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n595_), .A2(new_n597_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT16), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT76), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n582_), .A2(new_n583_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n616_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n622_), .B(KEYINPUT17), .Z(new_n629_));
  NAND2_X1  g428(.A1(new_n616_), .A2(new_n627_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT77), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n569_), .A2(new_n614_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n522_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n466_), .B(KEYINPUT103), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n481_), .A3(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT38), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n614_), .A2(new_n520_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n632_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n562_), .A2(new_n565_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT104), .B1(new_n477_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n473_), .A2(new_n475_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n471_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n279_), .ZN(new_n649_));
  AND4_X1   g448(.A1(new_n466_), .A2(new_n455_), .A3(new_n465_), .A4(new_n468_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n425_), .A2(new_n427_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n651_), .A2(new_n418_), .A3(new_n421_), .A4(new_n416_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n455_), .B1(new_n652_), .B2(new_n414_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n648_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656_));
  INV_X1    g455(.A(new_n644_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n643_), .B1(new_n645_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G1gat), .B1(new_n660_), .B2(new_n466_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n640_), .A2(new_n661_), .ZN(G1324gat));
  NAND2_X1  g461(.A1(new_n465_), .A2(new_n468_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n636_), .A2(new_n482_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n659_), .A2(new_n663_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(G8gat), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT39), .B(new_n482_), .C1(new_n659_), .C2(new_n663_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g469(.A1(new_n635_), .A2(G15gat), .A3(new_n649_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G15gat), .B1(new_n660_), .B2(new_n649_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(G1326gat));
  NAND3_X1  g475(.A1(new_n636_), .A2(new_n485_), .A3(new_n455_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n659_), .A2(new_n455_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(G22gat), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT42), .B(new_n485_), .C1(new_n659_), .C2(new_n455_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT105), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n633_), .A2(new_n644_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(new_n614_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n522_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n466_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n633_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(new_n614_), .A3(new_n520_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n655_), .B2(new_n569_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n692_), .B(new_n569_), .C1(new_n470_), .C2(new_n476_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT44), .B(new_n691_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n638_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n689_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(new_n663_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n686_), .A2(G36gat), .A3(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT45), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n698_), .A2(new_n663_), .A3(new_n699_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G36gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT46), .B(new_n705_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  NAND3_X1  g513(.A1(new_n700_), .A2(G43gat), .A3(new_n279_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n238_), .B1(new_n686_), .B2(new_n649_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT107), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g518(.A1(new_n686_), .A2(G50gat), .A3(new_n453_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n700_), .A2(new_n455_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n721_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT108), .B1(new_n721_), .B2(G50gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(G1331gat));
  NAND3_X1  g523(.A1(new_n690_), .A2(new_n614_), .A3(new_n521_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n645_), .B2(new_n658_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n466_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n655_), .A2(new_n520_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT109), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n569_), .A2(new_n633_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n614_), .A3(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n637_), .A2(G57gat), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n728_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT110), .Z(G1332gat));
  OR3_X1    g535(.A1(new_n732_), .A2(G64gat), .A3(new_n703_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n726_), .A2(new_n663_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G64gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT111), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n737_), .B(new_n744_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1333gat));
  OR3_X1    g545(.A1(new_n732_), .A2(G71gat), .A3(new_n649_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G71gat), .B1(new_n727_), .B2(new_n649_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  OR3_X1    g550(.A1(new_n732_), .A2(G78gat), .A3(new_n453_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G78gat), .B1(new_n727_), .B2(new_n453_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT50), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT50), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(G1335gat));
  AND4_X1   g555(.A1(new_n644_), .A2(new_n730_), .A3(new_n614_), .A4(new_n633_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n638_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n693_), .A2(new_n695_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n614_), .A2(new_n520_), .A3(new_n633_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n688_), .A2(G85gat), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT112), .Z(new_n763_));
  AOI21_X1  g562(.A(new_n758_), .B1(new_n761_), .B2(new_n763_), .ZN(G1336gat));
  INV_X1    g563(.A(G92gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n757_), .A2(new_n765_), .A3(new_n663_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n759_), .A2(new_n703_), .A3(new_n760_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(new_n767_), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n757_), .A2(new_n279_), .A3(new_n541_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n761_), .A2(new_n279_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n770_), .A2(KEYINPUT113), .A3(G99gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT113), .B1(new_n770_), .B2(G99gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT51), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n769_), .B(new_n775_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n757_), .A2(new_n542_), .A3(new_n455_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n761_), .A2(new_n455_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G106gat), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT52), .B(new_n542_), .C1(new_n761_), .C2(new_n455_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n778_), .B(new_n785_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n646_), .A2(new_n279_), .A3(new_n638_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n598_), .A2(new_n594_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(KEYINPUT55), .C1(new_n600_), .C2(new_n601_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n602_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n598_), .A2(new_n594_), .A3(new_n590_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n571_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n606_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .ZN(new_n799_));
  INV_X1    g598(.A(new_n498_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n506_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n505_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n509_), .B1(new_n497_), .B2(new_n800_), .ZN(new_n804_));
  OR3_X1    g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n508_), .A3(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(new_n609_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n602_), .A2(new_n793_), .B1(new_n571_), .B2(new_n795_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n607_), .B1(new_n809_), .B2(new_n792_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n799_), .A2(new_n808_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n799_), .A2(new_n808_), .A3(KEYINPUT58), .A4(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n569_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n798_), .A2(new_n819_), .A3(KEYINPUT56), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n811_), .B1(new_n810_), .B2(KEYINPUT115), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n520_), .A2(new_n609_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n611_), .A2(new_n807_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n657_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT118), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n644_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(KEYINPUT57), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n818_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n657_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n690_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n836_));
  INV_X1    g635(.A(new_n614_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n731_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n521_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n836_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n634_), .A2(new_n521_), .A3(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n788_), .B(new_n790_), .C1(new_n835_), .C2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n521_), .A2(new_n255_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n828_), .A2(new_n829_), .A3(KEYINPUT57), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n829_), .B1(new_n828_), .B2(KEYINPUT57), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n817_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n832_), .A2(new_n849_), .A3(new_n833_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT117), .B1(new_n828_), .B2(KEYINPUT57), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n632_), .B1(new_n848_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n840_), .A2(new_n842_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n789_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n844_), .B(new_n845_), .C1(new_n855_), .C2(new_n788_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n520_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n850_), .A2(new_n851_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n642_), .B1(new_n858_), .B2(new_n831_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n857_), .B(new_n790_), .C1(new_n859_), .C2(new_n843_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n255_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT119), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n856_), .A2(new_n864_), .A3(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1340gat));
  OAI21_X1  g665(.A(new_n257_), .B1(new_n837_), .B2(KEYINPUT60), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n855_), .B(new_n867_), .C1(KEYINPUT60), .C2(new_n257_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n858_), .A2(new_n831_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n843_), .B1(new_n869_), .B2(new_n632_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT59), .B1(new_n870_), .B2(new_n789_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n614_), .A3(new_n844_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n868_), .B1(new_n873_), .B2(new_n257_), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n855_), .A2(new_n249_), .A3(new_n690_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(new_n642_), .A3(new_n844_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n249_), .ZN(G1342gat));
  AOI21_X1  g677(.A(G134gat), .B1(new_n855_), .B2(new_n644_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n871_), .A2(new_n844_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n569_), .A2(G134gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT120), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n879_), .B1(new_n880_), .B2(new_n882_), .ZN(G1343gat));
  XNOR2_X1  g682(.A(KEYINPUT122), .B(G141gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n279_), .A2(new_n453_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n638_), .A2(new_n703_), .A3(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT121), .B1(new_n870_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n853_), .A2(new_n854_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889_));
  INV_X1    g688(.A(new_n886_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n884_), .B1(new_n892_), .B2(new_n857_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n884_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n520_), .B(new_n894_), .C1(new_n887_), .C2(new_n891_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1344gat));
  XNOR2_X1  g695(.A(KEYINPUT123), .B(G148gat), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n889_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n899_));
  AOI211_X1 g698(.A(KEYINPUT121), .B(new_n886_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n898_), .B1(new_n901_), .B2(new_n837_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n892_), .A2(new_n614_), .A3(new_n897_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1345gat));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n901_), .B2(new_n633_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n905_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n892_), .A2(new_n690_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1346gat));
  INV_X1    g708(.A(new_n569_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G162gat), .B1(new_n901_), .B2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n892_), .A2(new_n379_), .A3(new_n644_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1347gat));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n638_), .A2(new_n703_), .A3(new_n649_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n455_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n831_), .A2(new_n834_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n633_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n920_), .B2(new_n854_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n857_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n914_), .B1(new_n922_), .B2(G169gat), .ZN(new_n923_));
  AOI211_X1 g722(.A(KEYINPUT62), .B(new_n207_), .C1(new_n921_), .C2(new_n857_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n921_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT22), .B(G169gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n857_), .A2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT124), .ZN(new_n928_));
  OAI22_X1  g727(.A1(new_n923_), .A2(new_n924_), .B1(new_n925_), .B2(new_n928_), .ZN(G1348gat));
  AOI21_X1  g728(.A(G176gat), .B1(new_n921_), .B2(new_n614_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n870_), .A2(new_n455_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n916_), .A2(new_n208_), .A3(new_n837_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  NOR3_X1   g732(.A1(new_n925_), .A2(new_n323_), .A3(new_n632_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n931_), .A2(new_n690_), .A3(new_n915_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n226_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n921_), .A2(new_n213_), .A3(new_n644_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n921_), .A2(new_n569_), .ZN(new_n939_));
  AOI21_X1  g738(.A(KEYINPUT125), .B1(new_n939_), .B2(G190gat), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  INV_X1    g740(.A(G190gat), .ZN(new_n942_));
  AOI211_X1 g741(.A(new_n941_), .B(new_n942_), .C1(new_n921_), .C2(new_n569_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n938_), .B1(new_n940_), .B2(new_n943_), .ZN(G1351gat));
  NAND3_X1  g743(.A1(new_n885_), .A2(new_n466_), .A3(new_n663_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n870_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n857_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n614_), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT126), .B(G204gat), .Z(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(G1353gat));
  AOI211_X1 g750(.A(KEYINPUT63), .B(G211gat), .C1(new_n946_), .C2(new_n642_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(KEYINPUT63), .B(G211gat), .ZN(new_n953_));
  NOR4_X1   g752(.A1(new_n870_), .A2(new_n632_), .A3(new_n945_), .A4(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n952_), .A2(new_n954_), .ZN(G1354gat));
  AOI21_X1  g754(.A(G218gat), .B1(new_n946_), .B2(new_n644_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n569_), .A2(G218gat), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(KEYINPUT127), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n956_), .B1(new_n946_), .B2(new_n958_), .ZN(G1355gat));
endmodule


