//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OAI211_X1 g005(.A(KEYINPUT71), .B(KEYINPUT14), .C1(new_n202_), .C2(new_n203_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT72), .ZN(new_n210_));
  XOR2_X1   g009(.A(G1gat), .B(G8gat), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n215_));
  XOR2_X1   g014(.A(G71gat), .B(G78gat), .Z(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n215_), .A2(new_n216_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n212_), .B(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223_));
  XOR2_X1   g022(.A(G127gat), .B(G155gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G183gat), .B(G211gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n222_), .A2(new_n223_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(KEYINPUT17), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n222_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT83), .B(G113gat), .ZN(new_n234_));
  INV_X1    g033(.A(G120gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT84), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT84), .ZN(new_n243_));
  OR3_X1    g042(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n245_));
  INV_X1    g044(.A(G141gat), .ZN(new_n246_));
  INV_X1    g045(.A(G148gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n244_), .A2(new_n248_), .A3(new_n249_), .A4(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n242_), .A2(new_n243_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n241_), .A2(new_n253_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n239_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n238_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(KEYINPUT85), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n252_), .B2(new_n256_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n238_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(new_n262_), .A3(KEYINPUT4), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n264_), .B(new_n238_), .C1(new_n259_), .C2(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT94), .Z(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT95), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n258_), .A2(new_n262_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n267_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n263_), .A2(new_n265_), .A3(KEYINPUT95), .A4(new_n267_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G1gat), .B(G29gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(G57gat), .B(G85gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n270_), .A2(new_n273_), .A3(new_n274_), .A4(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G226gat), .A2(G233gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT92), .Z(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT19), .Z(new_n289_));
  NOR2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT79), .ZN(new_n291_));
  INV_X1    g090(.A(G169gat), .ZN(new_n292_));
  INV_X1    g091(.A(G176gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n291_), .B(KEYINPUT24), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT23), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT26), .B(G190gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT78), .B(G183gat), .Z(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT25), .ZN(new_n300_));
  NOR2_X1   g099(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n298_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n297_), .B(new_n302_), .C1(KEYINPUT24), .C2(new_n291_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n296_), .B1(G190gat), .B2(new_n299_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n293_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT22), .ZN(new_n307_));
  AOI21_X1  g106(.A(G176gat), .B1(new_n307_), .B2(KEYINPUT80), .ZN(new_n308_));
  OAI221_X1 g107(.A(new_n304_), .B1(KEYINPUT80), .B2(new_n306_), .C1(new_n292_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT21), .B1(new_n311_), .B2(KEYINPUT89), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n312_), .B(new_n314_), .C1(KEYINPUT21), .C2(new_n311_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT20), .B1(new_n310_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT25), .B(G183gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT93), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n298_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n290_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n323_), .B(new_n297_), .C1(KEYINPUT24), .C2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n296_), .B1(G183gat), .B2(G190gat), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n326_), .B(new_n306_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n319_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n289_), .B1(new_n318_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT20), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n310_), .B2(new_n317_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n289_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(new_n319_), .A3(new_n327_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT18), .B(G64gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G92gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n286_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n318_), .A2(new_n289_), .A3(new_n328_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n332_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n340_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n346_), .B(KEYINPUT27), .C1(new_n340_), .C2(new_n335_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G233gat), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n349_), .A2(KEYINPUT88), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(KEYINPUT88), .ZN(new_n351_));
  OAI21_X1  g150(.A(G228gat), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n259_), .A2(new_n261_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n317_), .B(new_n352_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n352_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n354_), .B1(new_n252_), .B2(new_n256_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(new_n319_), .B2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT90), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT91), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n359_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n353_), .A2(new_n354_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G22gat), .B(G50gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n368_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT87), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT87), .B1(new_n369_), .B2(new_n370_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n363_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G15gat), .B(G43gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G71gat), .B(G99gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n310_), .A2(KEYINPUT30), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n310_), .A2(KEYINPUT30), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT81), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n382_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(new_n381_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n376_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n388_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n381_), .B1(new_n393_), .B2(new_n390_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n391_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n376_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n359_), .A2(new_n361_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n362_), .B2(new_n359_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n373_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n398_), .B1(new_n373_), .B2(new_n401_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n285_), .B(new_n348_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n339_), .A2(KEYINPUT32), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n335_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n405_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n284_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT98), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT97), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  OR3_X1    g211(.A1(new_n283_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n282_), .B1(new_n271_), .B2(new_n267_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n263_), .A2(new_n272_), .A3(new_n265_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n341_), .A2(new_n342_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n283_), .A2(new_n412_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n283_), .B2(new_n412_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n413_), .A2(new_n417_), .A3(new_n418_), .A4(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n284_), .A2(new_n407_), .A3(KEYINPUT98), .A4(new_n406_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n410_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n398_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n373_), .A2(new_n401_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n233_), .B1(new_n404_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(G106gat), .ZN(new_n427_));
  INV_X1    g226(.A(G99gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT10), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G99gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT64), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n427_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT65), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT9), .ZN(new_n437_));
  INV_X1    g236(.A(G85gat), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n438_), .A2(G92gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(G92gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(KEYINPUT66), .A3(G92gat), .ZN(new_n442_));
  OR2_X1    g241(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n438_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n428_), .B2(new_n427_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n441_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT65), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n450_), .B(new_n427_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n436_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT67), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n436_), .A2(new_n454_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n439_), .A2(new_n440_), .ZN(new_n457_));
  OR3_X1    g256(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n457_), .B1(new_n460_), .B2(new_n448_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT8), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n456_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n219_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n463_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n219_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(KEYINPUT12), .A3(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n468_), .A2(KEYINPUT12), .A3(new_n219_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G230gat), .A2(G233gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n219_), .B1(new_n456_), .B2(new_n464_), .ZN(new_n476_));
  AOI211_X1 g275(.A(new_n466_), .B(new_n463_), .C1(new_n453_), .C2(new_n455_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n475_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G120gat), .B(G148gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G204gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT5), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(G176gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n483_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT13), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(new_n488_), .A3(new_n485_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G169gat), .B(G197gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G141gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT76), .ZN(new_n493_));
  INV_X1    g292(.A(G113gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(KEYINPUT75), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n210_), .B(new_n211_), .Z(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  INV_X1    g298(.A(G43gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G50gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n501_), .B(G50gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n212_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n497_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT74), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n503_), .B(KEYINPUT69), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT15), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n505_), .B(KEYINPUT69), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n513_), .A3(new_n212_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n497_), .A3(new_n504_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n496_), .B1(new_n508_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n504_), .A2(new_n506_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n497_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT74), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT74), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(new_n521_), .A3(new_n518_), .ZN(new_n522_));
  AND4_X1   g321(.A1(new_n496_), .A2(new_n520_), .A3(new_n515_), .A4(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n490_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n510_), .A2(new_n513_), .A3(new_n465_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT34), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT68), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n468_), .B2(new_n503_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n527_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n532_), .B1(new_n527_), .B2(new_n534_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT70), .B(G190gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G218gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT36), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n538_), .A2(new_n544_), .ZN(new_n545_));
  NOR4_X1   g344(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT36), .A4(new_n542_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT100), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n542_), .A2(KEYINPUT36), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n538_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT100), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n549_), .B(new_n550_), .C1(new_n538_), .C2(new_n544_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n426_), .A2(new_n526_), .A3(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(G1gat), .B1(new_n553_), .B2(new_n285_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT101), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT37), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n549_), .B(KEYINPUT37), .C1(new_n538_), .C2(new_n544_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n426_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n524_), .A2(KEYINPUT77), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n561_), .A2(new_n490_), .A3(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(new_n202_), .A3(new_n284_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT102), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n568_), .A2(KEYINPUT102), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n567_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n555_), .B(new_n571_), .C1(new_n569_), .C2(new_n567_), .ZN(G1324gat));
  OR2_X1    g371(.A1(new_n553_), .A2(new_n348_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT104), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT104), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(G8gat), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT39), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n348_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n566_), .A2(new_n203_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT103), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n574_), .A2(KEYINPUT39), .A3(G8gat), .A4(new_n575_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT40), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n578_), .A2(new_n581_), .A3(KEYINPUT40), .A4(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(G1325gat));
  OAI21_X1  g386(.A(G15gat), .B1(new_n553_), .B2(new_n423_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT105), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT41), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n566_), .A2(new_n398_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n591_), .B(new_n592_), .C1(G15gat), .C2(new_n593_), .ZN(G1326gat));
  OAI21_X1  g393(.A(G22gat), .B1(new_n553_), .B2(new_n424_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT106), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT42), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n597_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n424_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n566_), .A2(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n598_), .B(new_n599_), .C1(G22gat), .C2(new_n601_), .ZN(G1327gat));
  AOI21_X1  g401(.A(new_n552_), .B1(new_n404_), .B2(new_n425_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n490_), .A2(new_n565_), .A3(new_n232_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n606_), .A2(G29gat), .A3(new_n285_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n404_), .A2(new_n425_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n559_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT43), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT43), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n611_), .A3(new_n559_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT44), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT107), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n613_), .A2(new_n233_), .A3(new_n526_), .A4(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n611_), .B1(new_n608_), .B2(new_n559_), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT43), .B(new_n560_), .C1(new_n404_), .C2(new_n425_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n233_), .B(new_n526_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n284_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n607_), .B1(new_n623_), .B2(G29gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT108), .ZN(G1328gat));
  NOR3_X1   g424(.A1(new_n606_), .A2(G36gat), .A3(new_n348_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT45), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n616_), .A2(new_n621_), .A3(new_n579_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT109), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n628_), .A2(new_n629_), .A3(G36gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n628_), .B2(G36gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT46), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n627_), .B(KEYINPUT46), .C1(new_n630_), .C2(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1329gat));
  NOR3_X1   g435(.A1(new_n606_), .A2(G43gat), .A3(new_n423_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n622_), .A2(new_n398_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(G43gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g439(.A1(new_n622_), .A2(G50gat), .A3(new_n600_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n502_), .B1(new_n606_), .B2(new_n424_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1331gat));
  AND2_X1   g442(.A1(new_n426_), .A2(new_n560_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n490_), .A2(new_n525_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(G57gat), .B1(new_n648_), .B2(new_n284_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n233_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n608_), .A2(new_n490_), .A3(new_n552_), .A4(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n285_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n649_), .B1(G57gat), .B2(new_n652_), .ZN(G1332gat));
  OAI21_X1  g452(.A(G64gat), .B1(new_n651_), .B2(new_n348_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT48), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n348_), .A2(G64gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n647_), .B2(new_n656_), .ZN(G1333gat));
  OAI21_X1  g456(.A(G71gat), .B1(new_n651_), .B2(new_n423_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT110), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT49), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n648_), .A2(new_n398_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n661_), .B(new_n662_), .C1(G71gat), .C2(new_n663_), .ZN(G1334gat));
  OAI21_X1  g463(.A(G78gat), .B1(new_n651_), .B2(new_n424_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT50), .ZN(new_n666_));
  INV_X1    g465(.A(G78gat), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n645_), .A2(new_n424_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n644_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(G1335gat));
  NOR2_X1   g469(.A1(new_n645_), .A2(new_n232_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n603_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G85gat), .B1(new_n672_), .B2(new_n284_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT111), .Z(new_n674_));
  OR2_X1    g473(.A1(new_n613_), .A2(KEYINPUT112), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n613_), .A2(KEYINPUT112), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(new_n671_), .A3(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n285_), .A2(new_n438_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1336gat));
  AOI21_X1  g478(.A(G92gat), .B1(new_n672_), .B2(new_n579_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n348_), .B1(new_n443_), .B2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n677_), .B2(new_n682_), .ZN(G1337gat));
  NAND4_X1  g482(.A1(new_n675_), .A2(new_n398_), .A3(new_n671_), .A4(new_n676_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n433_), .A2(new_n434_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n423_), .A2(new_n685_), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n684_), .A2(G99gat), .B1(new_n672_), .B2(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n687_), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n688_));
  NOR2_X1   g487(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n689_));
  AND2_X1   g488(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n687_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n688_), .A2(new_n691_), .ZN(G1338gat));
  NAND3_X1  g491(.A1(new_n672_), .A2(new_n427_), .A3(new_n600_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n613_), .A2(new_n233_), .A3(new_n668_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT52), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(G106gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n694_), .B2(G106gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g498(.A(KEYINPUT114), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n487_), .A2(new_n489_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n650_), .A3(new_n560_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n702_), .B2(KEYINPUT54), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n559_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT54), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n704_), .A2(KEYINPUT114), .A3(new_n705_), .A4(new_n650_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(KEYINPUT54), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n703_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n497_), .B1(new_n514_), .B2(new_n504_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n517_), .A2(new_n518_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n495_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n520_), .A2(new_n515_), .A3(new_n522_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(new_n495_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT55), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n471_), .B1(new_n478_), .B2(KEYINPUT12), .ZN(new_n716_));
  INV_X1    g515(.A(new_n474_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT115), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT115), .B(new_n717_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT115), .B1(new_n716_), .B2(new_n717_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n470_), .A2(new_n717_), .A3(new_n472_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT55), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n473_), .A2(new_n719_), .A3(new_n474_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n722_), .A2(new_n483_), .A3(new_n727_), .A4(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n524_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n479_), .A2(new_n483_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n722_), .A2(new_n483_), .A3(new_n727_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n728_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n714_), .B1(new_n730_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n552_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT117), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n732_), .A2(new_n733_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n738_), .A2(new_n484_), .A3(new_n524_), .A4(new_n729_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n714_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n552_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n713_), .B1(new_n732_), .B2(KEYINPUT56), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n722_), .A2(new_n747_), .A3(new_n727_), .A4(new_n483_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n484_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT58), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n746_), .A2(KEYINPUT58), .A3(new_n484_), .A4(new_n748_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n559_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT118), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n741_), .A2(KEYINPUT57), .A3(new_n552_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT118), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n751_), .A2(new_n756_), .A3(new_n559_), .A4(new_n752_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n745_), .A2(new_n754_), .A3(new_n755_), .A4(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n708_), .B1(new_n758_), .B2(new_n233_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n579_), .A2(new_n285_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n402_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT59), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n565_), .A2(new_n494_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n745_), .A2(new_n753_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n745_), .A2(KEYINPUT119), .A3(new_n753_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n755_), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n708_), .B1(new_n768_), .B2(new_n233_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n761_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT59), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n762_), .B(new_n763_), .C1(new_n769_), .C2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n759_), .A2(new_n761_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n524_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n494_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n776_), .A3(KEYINPUT120), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1340gat));
  NAND2_X1  g580(.A1(new_n767_), .A2(new_n755_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT119), .B1(new_n745_), .B2(new_n753_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n233_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n708_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n771_), .A3(new_n770_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n490_), .A3(new_n762_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G120gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n235_), .B1(new_n701_), .B2(KEYINPUT60), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n774_), .B(new_n790_), .C1(KEYINPUT60), .C2(new_n235_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1341gat));
  AOI21_X1  g591(.A(G127gat), .B1(new_n774_), .B2(new_n232_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n787_), .A2(new_n762_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n232_), .A2(G127gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(G1342gat));
  AOI21_X1  g595(.A(G134gat), .B1(new_n774_), .B2(new_n736_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n559_), .A2(G134gat), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT121), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n794_), .B2(new_n799_), .ZN(G1343gat));
  INV_X1    g599(.A(new_n403_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n759_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT122), .B1(new_n802_), .B2(new_n760_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n804_));
  INV_X1    g603(.A(new_n760_), .ZN(new_n805_));
  NOR4_X1   g604(.A1(new_n759_), .A2(new_n804_), .A3(new_n801_), .A4(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n524_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G141gat), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n246_), .B(new_n524_), .C1(new_n803_), .C2(new_n806_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1344gat));
  OAI21_X1  g609(.A(new_n490_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G148gat), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n247_), .B(new_n490_), .C1(new_n803_), .C2(new_n806_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1345gat));
  OAI21_X1  g613(.A(new_n232_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT61), .B(G155gat), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT123), .Z(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n817_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n232_), .B(new_n819_), .C1(new_n803_), .C2(new_n806_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1346gat));
  OR2_X1    g620(.A1(new_n803_), .A2(new_n806_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n559_), .A2(G162gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT124), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n736_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n825_));
  INV_X1    g624(.A(G162gat), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n822_), .A2(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(G1347gat));
  NOR2_X1   g626(.A1(new_n348_), .A2(new_n284_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n786_), .A2(new_n524_), .A3(new_n402_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G169gat), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n786_), .A2(new_n402_), .A3(new_n828_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n524_), .A3(new_n305_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n829_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n835_), .A3(new_n836_), .ZN(G1348gat));
  OAI21_X1  g636(.A(new_n293_), .B1(new_n833_), .B2(new_n701_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n759_), .A2(new_n600_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n828_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n423_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n839_), .A2(G176gat), .A3(new_n490_), .A4(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n838_), .A2(new_n842_), .ZN(G1349gat));
  NOR3_X1   g642(.A1(new_n840_), .A2(new_n233_), .A3(new_n423_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n299_), .B1(new_n839_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n233_), .A2(new_n322_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n834_), .B2(new_n846_), .ZN(G1350gat));
  OAI21_X1  g646(.A(G190gat), .B1(new_n833_), .B2(new_n560_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n736_), .A2(new_n298_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n833_), .B2(new_n849_), .ZN(G1351gat));
  NOR3_X1   g649(.A1(new_n759_), .A2(new_n801_), .A3(new_n840_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n524_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n490_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT126), .Z(new_n856_));
  XOR2_X1   g655(.A(new_n854_), .B(new_n856_), .Z(G1353gat));
  NOR4_X1   g656(.A1(new_n759_), .A2(new_n233_), .A3(new_n801_), .A4(new_n840_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n859_));
  INV_X1    g658(.A(G211gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n860_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n858_), .A2(new_n861_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT127), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT127), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n858_), .A2(new_n866_), .A3(new_n861_), .A4(new_n863_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n858_), .A2(new_n861_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(G1354gat));
  AOI21_X1  g668(.A(G218gat), .B1(new_n851_), .B2(new_n736_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n851_), .A2(new_n559_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(G218gat), .B2(new_n871_), .ZN(G1355gat));
endmodule


