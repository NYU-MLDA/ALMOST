//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_;
  XOR2_X1   g000(.A(KEYINPUT82), .B(G176gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT23), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n207_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT26), .B(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G169gat), .B2(G176gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n217_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n212_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT81), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n210_), .A2(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(KEYINPUT81), .B(KEYINPUT23), .C1(new_n208_), .C2(new_n209_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OAI22_X1  g026(.A1(new_n206_), .A2(new_n213_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT30), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G15gat), .B(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  INV_X1    g033(.A(G71gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n232_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n231_), .B(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n236_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n243_), .A2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n242_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n243_), .A2(new_n244_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT85), .A3(new_n245_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT31), .Z(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(G99gat), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n238_), .A2(new_n241_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n205_), .B(new_n204_), .C1(new_n227_), .C2(new_n207_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n205_), .A2(KEYINPUT24), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n220_), .B1(new_n258_), .B2(KEYINPUT91), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT91), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n218_), .A2(new_n260_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n259_), .A2(new_n261_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT92), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n210_), .A2(new_n212_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(new_n262_), .B2(KEYINPUT92), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n257_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G197gat), .A2(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G197gat), .A2(G204gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT21), .A3(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G211gat), .B(G218gat), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  INV_X1    g073(.A(new_n270_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n274_), .B1(new_n275_), .B2(new_n268_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n276_), .A3(new_n272_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n267_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n278_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT19), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT96), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT96), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n279_), .A2(new_n281_), .A3(new_n287_), .A4(new_n284_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT20), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n228_), .B2(new_n278_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n267_), .B2(new_n278_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n283_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n288_), .A3(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G8gat), .B(G36gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT18), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n278_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT92), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n259_), .A2(new_n261_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n216_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n305_), .B2(new_n257_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n283_), .B1(new_n306_), .B2(new_n280_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n290_), .B(new_n284_), .C1(new_n267_), .C2(new_n278_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n307_), .A2(new_n297_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n298_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(new_n297_), .A3(new_n308_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n299_), .A2(new_n311_), .B1(new_n315_), .B2(new_n310_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT89), .ZN(new_n317_));
  XOR2_X1   g116(.A(G22gat), .B(G50gat), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(KEYINPUT1), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(KEYINPUT86), .A3(G155gat), .A4(G162gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(KEYINPUT1), .ZN(new_n325_));
  OR2_X1    g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n322_), .A2(new_n324_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G141gat), .B(G148gat), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330_));
  INV_X1    g129(.A(G141gat), .ZN(new_n331_));
  INV_X1    g130(.A(G148gat), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .A4(KEYINPUT87), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n334_));
  OAI22_X1  g133(.A1(new_n334_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n333_), .A2(new_n335_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n326_), .A2(new_n321_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n329_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT28), .B1(new_n343_), .B2(KEYINPUT29), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT88), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n327_), .A2(new_n328_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n344_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n345_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n319_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n344_), .A2(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT88), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n344_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n318_), .A3(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n346_), .A2(new_n348_), .ZN(new_n358_));
  OAI21_X1  g157(.A(G106gat), .B1(new_n358_), .B2(new_n300_), .ZN(new_n359_));
  INV_X1    g158(.A(G106gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n278_), .C1(new_n346_), .C2(new_n348_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n363_), .B(G78gat), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n359_), .A2(new_n364_), .A3(new_n361_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n317_), .B1(new_n357_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n352_), .A2(new_n356_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n371_), .A2(new_n368_), .A3(KEYINPUT89), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n371_), .A2(KEYINPUT90), .A3(new_n368_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT90), .B1(new_n371_), .B2(new_n368_), .ZN(new_n374_));
  OAI22_X1  g173(.A1(new_n370_), .A2(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n248_), .A2(new_n343_), .A3(new_n250_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n346_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n248_), .A2(new_n343_), .A3(new_n381_), .A4(new_n250_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT94), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n376_), .A2(new_n377_), .A3(KEYINPUT4), .ZN(new_n385_));
  INV_X1    g184(.A(new_n379_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n380_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT95), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n393_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n380_), .B(new_n395_), .C1(new_n384_), .C2(new_n387_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n316_), .A2(new_n375_), .A3(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n297_), .A2(KEYINPUT32), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n293_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(new_n397_), .C1(new_n400_), .C2(new_n312_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n297_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n309_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n313_), .A2(KEYINPUT93), .A3(new_n314_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n396_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n376_), .A2(new_n377_), .A3(new_n386_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n393_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n382_), .B(KEYINPUT94), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n385_), .A2(new_n379_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n396_), .B2(new_n407_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n405_), .A2(new_n406_), .A3(new_n408_), .A4(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n375_), .B1(new_n402_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n399_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI211_X1 g217(.A(KEYINPUT97), .B(new_n375_), .C1(new_n402_), .C2(new_n415_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n256_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT98), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n238_), .A2(new_n241_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n253_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n238_), .A2(new_n241_), .A3(new_n253_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n375_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n398_), .A3(new_n427_), .A4(new_n316_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT98), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n256_), .B(new_n429_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n421_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G43gat), .B(G50gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G36gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G29gat), .ZN(new_n436_));
  INV_X1    g235(.A(G29gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G36gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n434_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n437_), .A2(G36gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n435_), .A2(G29gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT73), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n433_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(KEYINPUT80), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G15gat), .B(G22gat), .ZN(new_n450_));
  INV_X1    g249(.A(G1gat), .ZN(new_n451_));
  INV_X1    g250(.A(G8gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT14), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G1gat), .B(G8gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n442_), .A2(KEYINPUT80), .A3(new_n447_), .ZN(new_n458_));
  OR3_X1    g257(.A1(new_n449_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n457_), .B1(new_n449_), .B2(new_n458_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G229gat), .A2(G233gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G141gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G169gat), .B(G197gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n442_), .A2(new_n447_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT15), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n456_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n460_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n464_), .B(new_n467_), .C1(new_n463_), .C2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n467_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n472_), .A2(new_n463_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n462_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n432_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G232gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT34), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT65), .ZN(new_n492_));
  OR2_X1    g291(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n360_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n491_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n493_), .A2(KEYINPUT65), .A3(new_n360_), .A4(new_n494_), .ZN(new_n497_));
  INV_X1    g296(.A(G85gat), .ZN(new_n498_));
  INV_X1    g297(.A(G92gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(KEYINPUT9), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G92gat), .ZN(new_n505_));
  OR2_X1    g304(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n503_), .A2(new_n508_), .A3(KEYINPUT67), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT67), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT66), .B(G85gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n505_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n513_), .B2(new_n502_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n496_), .B(new_n497_), .C1(new_n509_), .C2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n490_), .A2(KEYINPUT69), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT69), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n487_), .A2(new_n489_), .A3(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520_));
  AND2_X1   g319(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n521_));
  NOR2_X1   g320(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI22_X1  g322(.A1(KEYINPUT68), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n517_), .A2(new_n519_), .A3(new_n523_), .A4(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n500_), .A2(new_n501_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n516_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n524_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(new_n491_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n516_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n515_), .B1(new_n528_), .B2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n470_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n515_), .B(new_n448_), .C1(new_n528_), .C2(new_n532_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT76), .B1(new_n483_), .B2(new_n484_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n485_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n470_), .A2(new_n533_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n485_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(KEYINPUT75), .A3(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G190gat), .B(G218gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT74), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n538_), .A2(KEYINPUT75), .A3(new_n541_), .A4(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT77), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT37), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n456_), .B(new_n558_), .Z(new_n559_));
  AND2_X1   g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n563_), .B2(KEYINPUT11), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT70), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n563_), .B2(KEYINPUT11), .ZN(new_n566_));
  INV_X1    g365(.A(G64gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G57gat), .ZN(new_n568_));
  INV_X1    g367(.A(G57gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(G64gat), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n568_), .A2(new_n570_), .A3(new_n565_), .A4(KEYINPUT11), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n564_), .B1(new_n566_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n568_), .A2(new_n570_), .A3(KEYINPUT11), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT70), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n568_), .A2(new_n570_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT11), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n575_), .A2(new_n578_), .A3(new_n562_), .A4(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n559_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT78), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n581_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n580_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n573_), .A2(new_n579_), .A3(KEYINPUT71), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AOI211_X1 g393(.A(new_n587_), .B(new_n586_), .C1(new_n559_), .C2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n594_), .B2(new_n559_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n553_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(KEYINPUT77), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n557_), .A2(new_n597_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  INV_X1    g401(.A(new_n580_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n533_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT12), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT64), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n515_), .B(new_n580_), .C1(new_n528_), .C2(new_n532_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n533_), .A2(KEYINPUT12), .A3(new_n593_), .A4(new_n592_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n606_), .A2(new_n609_), .A3(new_n610_), .A4(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n604_), .A2(new_n610_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n608_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT5), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n612_), .A2(new_n614_), .A3(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n620_), .A2(KEYINPUT72), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT72), .B1(new_n620_), .B2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n602_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n622_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT72), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n620_), .A2(KEYINPUT72), .A3(new_n622_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(KEYINPUT13), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n601_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT79), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n480_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n451_), .A3(new_n397_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT38), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n631_), .A2(new_n479_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n597_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n555_), .B(KEYINPUT99), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n430_), .A2(new_n428_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n415_), .A2(new_n402_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT97), .B1(new_n646_), .B2(new_n375_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n416_), .A2(new_n417_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(new_n399_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n429_), .B1(new_n649_), .B2(new_n256_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n642_), .B(new_n644_), .C1(new_n645_), .C2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n642_), .B1(new_n431_), .B2(new_n644_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n641_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT101), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n641_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n655_), .A2(new_n397_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n637_), .B1(new_n658_), .B2(new_n451_), .ZN(G1324gat));
  INV_X1    g458(.A(new_n316_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n635_), .A2(new_n452_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(KEYINPUT39), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT102), .B1(new_n654_), .B2(new_n316_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n431_), .A2(new_n644_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT100), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n651_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n660_), .A4(new_n641_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n664_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n452_), .B1(new_n662_), .B2(KEYINPUT39), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n663_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n663_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n671_), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n673_), .B(new_n674_), .C1(new_n664_), .C2(new_n669_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n661_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT40), .B(new_n661_), .C1(new_n672_), .C2(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  OR3_X1    g479(.A1(new_n634_), .A2(G15gat), .A3(new_n256_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n655_), .A2(new_n426_), .A3(new_n657_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT41), .B1(new_n682_), .B2(G15gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT104), .B(new_n681_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1326gat));
  NAND3_X1  g488(.A1(new_n655_), .A2(new_n375_), .A3(new_n657_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n690_), .A2(new_n691_), .A3(G22gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n690_), .B2(G22gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n427_), .A2(G22gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT105), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n692_), .A2(new_n693_), .B1(new_n634_), .B2(new_n695_), .ZN(G1327gat));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n431_), .B1(KEYINPUT107), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n557_), .A2(new_n600_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n698_), .B(new_n699_), .C1(KEYINPUT107), .C2(new_n431_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n431_), .A2(new_n699_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n639_), .A2(new_n597_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n704_), .A4(new_n705_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n397_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G29gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n640_), .A2(new_n555_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(new_n631_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n480_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n437_), .A3(new_n397_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n711_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT108), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n711_), .A2(new_n719_), .A3(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1328gat));
  NAND3_X1  g520(.A1(new_n715_), .A2(new_n435_), .A3(new_n660_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT45), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n708_), .A2(new_n660_), .A3(new_n709_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G36gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n725_), .A3(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  NAND4_X1  g529(.A1(new_n708_), .A2(G43gat), .A3(new_n426_), .A4(new_n709_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n714_), .A2(new_n256_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(G43gat), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g533(.A(G50gat), .B1(new_n715_), .B2(new_n375_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n708_), .A2(new_n709_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n375_), .A2(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n631_), .A2(new_n479_), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n640_), .B(new_n739_), .C1(new_n666_), .C2(new_n651_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n398_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n432_), .A2(new_n478_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n631_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n601_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT109), .Z(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n569_), .A3(new_n397_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n742_), .A2(new_n749_), .ZN(G1332gat));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n567_), .A3(new_n660_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G64gat), .B1(new_n741_), .B2(new_n316_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT48), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(KEYINPUT48), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1333gat));
  NAND3_X1  g554(.A1(new_n748_), .A2(new_n235_), .A3(new_n426_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G71gat), .B1(new_n741_), .B2(new_n256_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(KEYINPUT49), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(KEYINPUT49), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n758_), .B2(new_n759_), .ZN(G1334gat));
  OR3_X1    g559(.A1(new_n747_), .A2(G78gat), .A3(new_n427_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G78gat), .B1(new_n741_), .B2(new_n427_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT50), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT50), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1335gat));
  AND2_X1   g564(.A1(new_n700_), .A2(new_n704_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n739_), .A2(new_n597_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n398_), .B(new_n768_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n744_), .A2(new_n712_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n743_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n397_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n769_), .A2(new_n773_), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n768_), .B2(new_n316_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n499_), .A3(new_n660_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n768_), .B2(new_n256_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n772_), .A2(new_n493_), .A3(new_n494_), .A4(new_n426_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g580(.A1(new_n772_), .A2(new_n360_), .A3(new_n375_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n700_), .A2(new_n375_), .A3(new_n704_), .A4(new_n767_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(G106gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(G106gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g587(.A1(new_n426_), .A2(new_n397_), .A3(new_n427_), .A4(new_n316_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n462_), .B1(new_n472_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n790_), .B2(new_n472_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n467_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n473_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n592_), .A2(KEYINPUT12), .A3(new_n593_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n495_), .A2(new_n492_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n490_), .A3(new_n497_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT67), .B1(new_n503_), .B2(new_n508_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n513_), .A2(new_n510_), .A3(new_n502_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n487_), .A2(new_n489_), .A3(new_n518_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n518_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n529_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT8), .B1(new_n806_), .B2(new_n526_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n530_), .A2(new_n531_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n803_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n610_), .B1(new_n798_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT12), .B1(new_n533_), .B2(new_n603_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n810_), .A2(new_n608_), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n608_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(KEYINPUT55), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  NOR4_X1   g614(.A1(new_n810_), .A2(new_n811_), .A3(new_n815_), .A4(new_n608_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n619_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n813_), .A2(KEYINPUT55), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n612_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n816_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n619_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n819_), .A2(new_n820_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n478_), .A2(new_n622_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n797_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT57), .A3(new_n599_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n824_), .B2(new_n619_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n827_), .B1(new_n833_), .B2(KEYINPUT110), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n819_), .A2(new_n825_), .A3(new_n820_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n796_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n836_), .B2(new_n555_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n794_), .A2(new_n473_), .A3(new_n622_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n818_), .B(new_n621_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT58), .B(new_n840_), .C1(new_n833_), .C2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n699_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n819_), .A2(new_n825_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT58), .B1(new_n844_), .B2(new_n840_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n839_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n840_), .B1(new_n833_), .B2(new_n841_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n849_), .A2(KEYINPUT112), .A3(new_n699_), .A4(new_n842_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n640_), .B1(new_n838_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n632_), .B2(new_n479_), .ZN(new_n854_));
  NOR4_X1   g653(.A1(new_n601_), .A2(new_n631_), .A3(KEYINPUT54), .A4(new_n478_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n789_), .B1(new_n852_), .B2(new_n857_), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT113), .Z(new_n859_));
  AOI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n478_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n831_), .A2(new_n837_), .A3(new_n846_), .A4(new_n850_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n856_), .B1(new_n864_), .B2(new_n640_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT114), .B(KEYINPUT59), .C1(new_n865_), .C2(new_n789_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n831_), .B(new_n837_), .C1(new_n845_), .C2(new_n843_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n856_), .B1(new_n868_), .B2(new_n640_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n869_), .A2(KEYINPUT59), .A3(new_n789_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n867_), .A2(KEYINPUT115), .A3(new_n871_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(G113gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n478_), .B2(KEYINPUT116), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(KEYINPUT116), .B2(new_n878_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n860_), .B1(new_n877_), .B2(new_n880_), .ZN(G1340gat));
  OAI21_X1  g680(.A(G120gat), .B1(new_n872_), .B2(new_n744_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n859_), .ZN(new_n883_));
  INV_X1    g682(.A(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n744_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(KEYINPUT60), .B2(new_n884_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n882_), .B1(new_n883_), .B2(new_n886_), .ZN(G1341gat));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT115), .B1(new_n867_), .B2(new_n871_), .ZN(new_n889_));
  AOI211_X1 g688(.A(new_n873_), .B(new_n870_), .C1(new_n863_), .C2(new_n866_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n597_), .A2(G127gat), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G127gat), .B1(new_n859_), .B2(new_n597_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n888_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n893_), .ZN(new_n895_));
  OAI211_X1 g694(.A(KEYINPUT117), .B(new_n895_), .C1(new_n876_), .C2(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1342gat));
  INV_X1    g696(.A(new_n699_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G134gat), .B1(new_n876_), .B2(new_n898_), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n883_), .A2(G134gat), .A3(new_n644_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1343gat));
  NAND3_X1  g700(.A1(new_n256_), .A2(new_n397_), .A3(new_n375_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n865_), .A2(new_n660_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n478_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT118), .B(G141gat), .Z(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1344gat));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n631_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT119), .B(G148gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1345gat));
  NAND2_X1  g708(.A1(new_n903_), .A2(new_n597_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT61), .B(G155gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1346gat));
  AOI21_X1  g711(.A(G162gat), .B1(new_n903_), .B2(new_n643_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n699_), .A2(G162gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT120), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n903_), .B2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT121), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n869_), .A2(new_n375_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n426_), .A2(new_n398_), .A3(new_n660_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n918_), .A2(new_n203_), .A3(new_n478_), .A4(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(G169gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n868_), .A2(new_n640_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n857_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n920_), .A2(new_n478_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT122), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n924_), .A2(new_n427_), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n922_), .B1(new_n927_), .B2(KEYINPUT123), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n918_), .A2(new_n926_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n928_), .A2(new_n929_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n929_), .B1(new_n928_), .B2(new_n932_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n921_), .B1(new_n933_), .B2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT124), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n937_), .B(new_n921_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1348gat));
  INV_X1    g738(.A(new_n918_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n919_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n631_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n865_), .A2(new_n375_), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n920_), .A2(G176gat), .A3(new_n631_), .ZN(new_n944_));
  AOI22_X1  g743(.A1(new_n942_), .A2(new_n202_), .B1(new_n943_), .B2(new_n944_), .ZN(G1349gat));
  NOR4_X1   g744(.A1(new_n940_), .A2(new_n214_), .A3(new_n640_), .A4(new_n919_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n946_), .A2(new_n947_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n919_), .A2(new_n640_), .ZN(new_n950_));
  AOI21_X1  g749(.A(G183gat), .B1(new_n943_), .B2(new_n950_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n948_), .A2(new_n949_), .A3(new_n951_), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n941_), .A2(new_n643_), .A3(new_n215_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n940_), .A2(new_n898_), .A3(new_n919_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n209_), .ZN(G1351gat));
  NAND4_X1  g754(.A1(new_n256_), .A2(new_n398_), .A3(new_n375_), .A4(new_n660_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n865_), .A2(new_n956_), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT126), .Z(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n478_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n631_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g761(.A1(new_n958_), .A2(new_n597_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  AND2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n963_), .A2(new_n964_), .A3(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n966_), .B1(new_n963_), .B2(new_n964_), .ZN(G1354gat));
  NAND2_X1  g766(.A1(new_n958_), .A2(new_n643_), .ZN(new_n968_));
  XOR2_X1   g767(.A(KEYINPUT127), .B(G218gat), .Z(new_n969_));
  NOR2_X1   g768(.A1(new_n898_), .A2(new_n969_), .ZN(new_n970_));
  AOI22_X1  g769(.A1(new_n968_), .A2(new_n969_), .B1(new_n958_), .B2(new_n970_), .ZN(G1355gat));
endmodule


