//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT7), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT66), .B(KEYINPUT6), .Z(new_n208_));
  OAI21_X1  g007(.A(new_n205_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n208_), .A2(new_n207_), .ZN(new_n210_));
  OAI211_X1 g009(.A(KEYINPUT8), .B(new_n203_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n202_), .B1(KEYINPUT9), .B2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G85gat), .Z(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(new_n212_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n206_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT10), .B(G99gat), .Z(new_n221_));
  AOI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G29gat), .B(G36gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n204_), .B(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n203_), .B1(new_n228_), .B2(new_n219_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n211_), .A2(new_n223_), .A3(new_n226_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G232gat), .A2(G233gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT34), .Z(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n211_), .A2(new_n223_), .A3(new_n231_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n226_), .B(KEYINPUT15), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  AOI211_X1 g040(.A(new_n234_), .B(new_n235_), .C1(new_n232_), .C2(KEYINPUT69), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G190gat), .B(G218gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G134gat), .B(G162gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(KEYINPUT36), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n242_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n243_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n246_), .B(KEYINPUT36), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT37), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT37), .B1(new_n253_), .B2(new_n254_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G57gat), .B(G64gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n259_));
  XOR2_X1   g058(.A(G71gat), .B(G78gat), .Z(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n260_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G231gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G8gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT71), .ZN(new_n268_));
  OR2_X1    g067(.A1(G15gat), .A2(G22gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G15gat), .A2(G22gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G1gat), .A2(G8gat), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n269_), .A2(new_n270_), .B1(KEYINPUT14), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n268_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n266_), .B(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G127gat), .B(G155gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G183gat), .B(G211gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT17), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n266_), .A2(new_n274_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n266_), .A2(new_n274_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n283_), .A2(KEYINPUT17), .A3(new_n280_), .A4(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n257_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n292_));
  AND2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT86), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(G141gat), .A3(G148gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G141gat), .ZN(new_n303_));
  INV_X1    g102(.A(G148gat), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n293_), .A2(KEYINPUT1), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n297_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n299_), .A2(new_n301_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(KEYINPUT2), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT87), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT3), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT87), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n312_), .B(new_n314_), .C1(G141gat), .C2(G148gat), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n311_), .A2(new_n303_), .A3(new_n304_), .A4(KEYINPUT3), .ZN(new_n316_));
  NAND3_X1  g115(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT89), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT89), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n315_), .A2(new_n316_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT2), .B1(new_n299_), .B2(new_n301_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT88), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n310_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n307_), .B1(new_n324_), .B2(new_n295_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n292_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n313_), .A2(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n311_), .A2(KEYINPUT3), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n316_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n318_), .A2(new_n320_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n330_), .B(new_n331_), .C1(new_n322_), .C2(KEYINPUT88), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n322_), .A2(KEYINPUT88), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n295_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  AND4_X1   g133(.A1(new_n292_), .A2(new_n334_), .A3(new_n326_), .A4(new_n306_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G22gat), .B(G50gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n327_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n306_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT28), .B1(new_n339_), .B2(KEYINPUT29), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n325_), .A2(new_n292_), .A3(new_n326_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT92), .B1(new_n338_), .B2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G78gat), .B(G106gat), .Z(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n337_), .B1(new_n327_), .B2(new_n335_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n341_), .A3(new_n336_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT92), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(G197gat), .A2(G204gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT21), .ZN(new_n353_));
  AND2_X1   g152(.A1(G197gat), .A2(G204gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n352_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT90), .ZN(new_n359_));
  INV_X1    g158(.A(G218gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G211gat), .ZN(new_n361_));
  INV_X1    g160(.A(G211gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(G218gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n364_), .A2(KEYINPUT21), .A3(new_n350_), .A4(new_n351_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n358_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n359_), .B1(new_n358_), .B2(new_n365_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(KEYINPUT29), .B2(new_n339_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT91), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n339_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n358_), .A2(new_n365_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n369_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n371_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n346_), .A2(new_n347_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n344_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(KEYINPUT92), .A3(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n345_), .A2(new_n349_), .A3(new_n378_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n349_), .A2(new_n378_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n379_), .B2(KEYINPUT92), .ZN(new_n384_));
  AOI211_X1 g183(.A(new_n348_), .B(new_n344_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT19), .Z(new_n393_));
  NOR2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT93), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(KEYINPUT24), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT24), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT93), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n394_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT25), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G183gat), .ZN(new_n401_));
  INV_X1    g200(.A(G190gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT26), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT26), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(G190gat), .ZN(new_n405_));
  INV_X1    g204(.A(G183gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT25), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n401_), .A2(new_n403_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G169gat), .ZN(new_n409_));
  INV_X1    g208(.A(G176gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n397_), .A2(KEYINPUT93), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n395_), .A2(KEYINPUT24), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .A4(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n399_), .A2(new_n408_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G183gat), .A2(G190gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(KEYINPUT23), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(KEYINPUT23), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(G183gat), .A3(G190gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n423_), .B2(new_n417_), .ZN(new_n424_));
  OR2_X1    g223(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n409_), .A2(KEYINPUT22), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT22), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G169gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n414_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n420_), .A2(new_n422_), .B1(new_n406_), .B2(new_n402_), .ZN(new_n432_));
  OAI22_X1  g231(.A1(new_n416_), .A2(new_n424_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT20), .B(new_n393_), .C1(new_n433_), .C2(new_n375_), .ZN(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT79), .B(G176gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT22), .B(G169gat), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n435_), .A2(new_n436_), .B1(G169gat), .B2(G176gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n438_), .A2(new_n439_), .A3(G190gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n437_), .B1(new_n424_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(KEYINPUT76), .A2(KEYINPUT77), .A3(G183gat), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n442_), .B(KEYINPUT25), .C1(KEYINPUT76), .C2(G183gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n400_), .A2(KEYINPUT77), .A3(G183gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT26), .B(G190gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n414_), .A2(KEYINPUT24), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(new_n394_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n420_), .A2(new_n422_), .B1(new_n397_), .B2(new_n394_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n411_), .A2(KEYINPUT78), .A3(KEYINPUT24), .A4(new_n414_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n441_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n434_), .B1(new_n453_), .B2(new_n368_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n441_), .B(new_n452_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n433_), .B2(new_n375_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n393_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n391_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n457_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n393_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n367_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n358_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n453_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n375_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n431_), .A2(new_n432_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n466_), .B(new_n467_), .C1(new_n424_), .C2(new_n416_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n465_), .A2(KEYINPUT20), .A3(new_n393_), .A4(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n391_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n459_), .A2(new_n471_), .A3(KEYINPUT94), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT94), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(new_n391_), .C1(new_n454_), .C2(new_n458_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G225gat), .A2(G233gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(G127gat), .B(G134gat), .Z(new_n477_));
  XOR2_X1   g276(.A(G113gat), .B(G120gat), .Z(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n325_), .B2(new_n480_), .ZN(new_n481_));
  AND4_X1   g280(.A1(new_n480_), .A2(new_n334_), .A3(new_n479_), .A4(new_n306_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n476_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G1gat), .B(G29gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G85gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT0), .B(G57gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(KEYINPUT4), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n334_), .A2(new_n480_), .A3(new_n306_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n479_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n325_), .A2(new_n480_), .A3(new_n479_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n339_), .A2(new_n488_), .A3(new_n479_), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n476_), .B(KEYINPUT96), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n483_), .B(new_n487_), .C1(new_n493_), .C2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT33), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT4), .B1(new_n481_), .B2(new_n482_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n494_), .A2(new_n495_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n502_), .A2(KEYINPUT33), .A3(new_n483_), .A4(new_n487_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n491_), .A2(new_n492_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n487_), .B1(new_n504_), .B2(new_n495_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n494_), .A2(new_n476_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n493_), .B2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n475_), .A2(new_n499_), .A3(new_n503_), .A4(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n391_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n462_), .A2(new_n469_), .A3(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n455_), .A2(new_n457_), .A3(new_n393_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT20), .B1(new_n433_), .B2(new_n375_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT97), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n433_), .C2(new_n375_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n465_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n513_), .B1(new_n518_), .B2(new_n461_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n512_), .B1(new_n519_), .B2(new_n511_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n487_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n493_), .A2(new_n496_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n483_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n521_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n520_), .B1(new_n524_), .B2(new_n497_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n508_), .B1(new_n525_), .B2(KEYINPUT98), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT98), .ZN(new_n527_));
  AOI211_X1 g326(.A(new_n527_), .B(new_n520_), .C1(new_n497_), .C2(new_n524_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n387_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n497_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n475_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n533_));
  NAND2_X1  g332(.A1(new_n518_), .A2(new_n461_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n513_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n470_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n471_), .A2(KEYINPUT27), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT99), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n514_), .A2(new_n515_), .B1(new_n368_), .B2(new_n453_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n393_), .B1(new_n539_), .B2(new_n517_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n391_), .B1(new_n540_), .B2(new_n513_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT99), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(KEYINPUT27), .A4(new_n471_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n532_), .A2(new_n533_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n531_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n529_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G43gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G227gat), .A2(G233gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(G71gat), .ZN(new_n550_));
  INV_X1    g349(.A(G71gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(G227gat), .A3(G233gat), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n550_), .A2(new_n552_), .A3(G99gat), .ZN(new_n553_));
  AOI21_X1  g352(.A(G99gat), .B1(new_n550_), .B2(new_n552_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n548_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n552_), .ZN(new_n556_));
  INV_X1    g355(.A(G99gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n550_), .A2(new_n552_), .A3(G99gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n547_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n441_), .A2(KEYINPUT30), .A3(new_n452_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT30), .B1(new_n441_), .B2(new_n452_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n453_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n441_), .A2(KEYINPUT30), .A3(new_n452_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n571_), .A2(new_n572_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT83), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n566_), .B1(new_n568_), .B2(new_n567_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n571_), .A2(new_n572_), .A3(new_n563_), .A4(new_n565_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT83), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n479_), .B(KEYINPUT31), .Z(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT84), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT85), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n575_), .A2(new_n576_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n581_), .B1(new_n587_), .B2(KEYINPUT83), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n583_), .A3(new_n578_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n585_), .A2(new_n586_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n586_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n530_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n538_), .A2(new_n543_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n472_), .A2(new_n474_), .A3(new_n533_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n595_), .A2(new_n382_), .A3(new_n386_), .A4(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT101), .B1(new_n594_), .B2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n588_), .A2(new_n578_), .B1(new_n583_), .B2(new_n582_), .ZN(new_n599_));
  AND4_X1   g398(.A1(new_n583_), .A2(new_n574_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT85), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n585_), .A2(new_n586_), .A3(new_n589_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n530_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n387_), .A4(new_n544_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n546_), .A2(new_n592_), .B1(new_n598_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n273_), .B(new_n226_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n274_), .A2(new_n239_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n273_), .A2(new_n226_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n608_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G113gat), .B(G141gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G169gat), .B(G197gat), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n614_), .B(new_n615_), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n610_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT75), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n610_), .A2(new_n613_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n616_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n620_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(KEYINPUT75), .A3(new_n617_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n606_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n264_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(new_n238_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n238_), .A2(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT12), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(KEYINPUT12), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n238_), .A2(new_n627_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n238_), .A2(new_n627_), .ZN(new_n636_));
  OAI211_X1 g435(.A(G230gat), .B(G233gat), .C1(new_n635_), .C2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT5), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n640_), .B(new_n641_), .Z(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT67), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n638_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT13), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n638_), .A2(new_n644_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n643_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n648_), .A2(new_n646_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n291_), .A2(new_n625_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT38), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n593_), .A2(G1gat), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n606_), .A2(new_n253_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n651_), .A2(new_n624_), .A3(new_n286_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n593_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n654_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT102), .ZN(G1324gat));
  INV_X1    g462(.A(new_n544_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n657_), .A2(new_n664_), .A3(new_n658_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G8gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT39), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n653_), .A2(G8gat), .A3(new_n544_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n659_), .B2(new_n592_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT41), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n653_), .A2(G15gat), .A3(new_n592_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  XOR2_X1   g473(.A(new_n387_), .B(KEYINPUT103), .Z(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n653_), .A2(G22gat), .A3(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n657_), .A2(new_n658_), .A3(new_n675_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n678_), .A2(G22gat), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n678_), .B2(G22gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT105), .ZN(G1327gat));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n606_), .B2(new_n257_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n255_), .A2(new_n256_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n598_), .A2(new_n605_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n592_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n529_), .B2(new_n545_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n685_), .B(new_n686_), .C1(new_n687_), .C2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n684_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n618_), .B(new_n622_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n286_), .B(KEYINPUT73), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n647_), .A2(new_n650_), .A3(new_n692_), .A4(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT106), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n691_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(KEYINPUT107), .A3(new_n530_), .A4(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n691_), .B2(new_n696_), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n698_), .B(new_n695_), .C1(new_n684_), .C2(new_n690_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT107), .B1(new_n705_), .B2(new_n530_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT108), .B1(new_n702_), .B2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n699_), .A2(new_n530_), .A3(new_n700_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(G29gat), .A4(new_n701_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n707_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n253_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n288_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT109), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n651_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n625_), .A2(new_n717_), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n718_), .A2(G29gat), .A3(new_n593_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n719_), .ZN(G1328gat));
  INV_X1    g519(.A(G36gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n705_), .B2(new_n664_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n718_), .A2(G36gat), .A3(new_n544_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT45), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  OR3_X1    g524(.A1(new_n722_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  NAND3_X1  g527(.A1(new_n705_), .A2(G43gat), .A3(new_n688_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n718_), .A2(new_n592_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(G43gat), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g531(.A(G50gat), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n387_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n625_), .A2(new_n717_), .A3(new_n675_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n705_), .A2(new_n734_), .B1(new_n735_), .B2(new_n733_), .ZN(G1331gat));
  NAND4_X1  g535(.A1(new_n657_), .A2(new_n624_), .A3(new_n651_), .A4(new_n288_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n593_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n291_), .A2(new_n651_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT110), .Z(new_n740_));
  NOR2_X1   g539(.A1(new_n606_), .A2(new_n692_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n593_), .A2(G57gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n738_), .B1(new_n742_), .B2(new_n743_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n737_), .B2(new_n544_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT48), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n544_), .A2(G64gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n742_), .B2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n737_), .B2(new_n592_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT49), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n688_), .A2(new_n551_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n742_), .B2(new_n751_), .ZN(G1334gat));
  OAI21_X1  g551(.A(G78gat), .B1(new_n737_), .B2(new_n676_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT50), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n676_), .A2(G78gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n742_), .B2(new_n755_), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n716_), .A2(new_n652_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n741_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n530_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n652_), .A2(new_n692_), .A3(new_n288_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n691_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n593_), .A2(new_n214_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(G1336gat));
  NAND2_X1  g564(.A1(new_n759_), .A2(new_n664_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n766_), .A2(KEYINPUT111), .A3(new_n212_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT111), .B1(new_n766_), .B2(new_n212_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n664_), .A2(G92gat), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n767_), .A2(new_n768_), .B1(new_n762_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT112), .ZN(G1337gat));
  AND2_X1   g570(.A1(new_n688_), .A2(new_n221_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT114), .B1(new_n759_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n763_), .A2(new_n688_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G99gat), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT113), .B(new_n557_), .C1(new_n763_), .C2(new_n688_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT51), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1338gat));
  INV_X1    g581(.A(new_n387_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n759_), .A2(new_n220_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n763_), .A2(new_n783_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(G106gat), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT52), .B(new_n220_), .C1(new_n763_), .C2(new_n783_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n784_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT115), .B1(new_n693_), .B2(new_n692_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n288_), .A2(new_n796_), .A3(new_n624_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n795_), .A2(new_n797_), .A3(new_n650_), .A4(new_n647_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n794_), .B1(new_n799_), .B2(new_n257_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n686_), .A2(new_n798_), .A3(KEYINPUT54), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n607_), .A2(new_n608_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n611_), .A2(new_n612_), .A3(new_n609_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n620_), .A3(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(new_n617_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n645_), .A2(KEYINPUT118), .A3(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT12), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n635_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n628_), .B1(new_n815_), .B2(new_n631_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n813_), .B1(new_n816_), .B2(KEYINPUT55), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n634_), .A2(KEYINPUT116), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(KEYINPUT55), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n630_), .B(new_n814_), .ZN(new_n821_));
  OAI211_X1 g620(.A(G230gat), .B(G233gat), .C1(new_n821_), .C2(new_n636_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n817_), .A2(new_n819_), .A3(new_n820_), .A4(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n642_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n642_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n825_), .A2(new_n826_), .A3(KEYINPUT117), .ZN(new_n827_));
  INV_X1    g626(.A(new_n642_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n634_), .A2(new_n637_), .A3(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n621_), .A2(new_n623_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n823_), .A2(new_n642_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n812_), .B1(new_n827_), .B2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT57), .A3(new_n714_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n834_), .A2(new_n835_), .A3(new_n824_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n830_), .B1(new_n826_), .B2(KEYINPUT117), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n811_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n839_), .B1(new_n842_), .B2(new_n253_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n806_), .A2(new_n829_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n806_), .A2(KEYINPUT119), .A3(new_n829_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT58), .B(new_n848_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n686_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n838_), .A2(new_n843_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n802_), .B1(new_n854_), .B2(new_n286_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n592_), .A2(new_n593_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n597_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(G113gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n692_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT59), .B1(new_n855_), .B2(new_n858_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT57), .B1(new_n837_), .B2(new_n714_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n851_), .A2(new_n686_), .A3(new_n852_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT120), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n843_), .A2(new_n867_), .A3(new_n853_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n838_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n802_), .B1(new_n869_), .B2(new_n693_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n858_), .A2(KEYINPUT59), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n692_), .B(new_n863_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n862_), .B1(new_n873_), .B2(new_n861_), .ZN(G1340gat));
  OAI21_X1  g673(.A(new_n863_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G120gat), .B1(new_n875_), .B2(new_n652_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n877_));
  AOI21_X1  g676(.A(G120gat), .B1(new_n651_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT121), .B1(new_n877_), .B2(G120gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n878_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n876_), .B1(new_n859_), .B2(new_n882_), .ZN(G1341gat));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n860_), .A2(new_n884_), .A3(new_n288_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n286_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n863_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n885_), .B1(new_n888_), .B2(new_n884_), .ZN(G1342gat));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n257_), .A2(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n863_), .B(new_n891_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n859_), .B2(new_n714_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT122), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n892_), .A2(new_n896_), .A3(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1343gat));
  NOR2_X1   g697(.A1(new_n688_), .A2(new_n387_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n544_), .A2(new_n530_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n855_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n692_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n651_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g705(.A1(new_n902_), .A2(new_n288_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT61), .B(G155gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1346gat));
  INV_X1    g708(.A(G162gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n902_), .A2(new_n910_), .A3(new_n253_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n855_), .A2(new_n257_), .A3(new_n900_), .A4(new_n901_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n910_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT123), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n911_), .B(new_n915_), .C1(new_n910_), .C2(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n544_), .A2(new_n530_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n688_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n675_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n870_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n692_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(G169gat), .A3(new_n925_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n870_), .A2(new_n624_), .A3(new_n921_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n436_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n924_), .B1(new_n927_), .B2(new_n409_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n926_), .A2(new_n928_), .A3(new_n929_), .ZN(G1348gat));
  NOR3_X1   g729(.A1(new_n855_), .A2(new_n783_), .A3(new_n919_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n652_), .A2(new_n410_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT125), .ZN(new_n934_));
  INV_X1    g733(.A(new_n435_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n922_), .B2(new_n651_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n934_), .A2(new_n936_), .ZN(G1349gat));
  AOI21_X1  g736(.A(new_n286_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n931_), .A2(new_n288_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n438_), .A2(new_n439_), .ZN(new_n940_));
  AOI22_X1  g739(.A1(new_n922_), .A2(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(G1350gat));
  NAND3_X1  g740(.A1(new_n922_), .A2(new_n445_), .A3(new_n253_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n870_), .A2(new_n257_), .A3(new_n921_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n402_), .ZN(G1351gat));
  XNOR2_X1  g743(.A(KEYINPUT127), .B(G197gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n854_), .A2(new_n286_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n802_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n948_), .A2(new_n899_), .A3(new_n918_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n900_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n952_), .A2(KEYINPUT126), .A3(new_n918_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n945_), .B1(new_n954_), .B2(new_n692_), .ZN(new_n955_));
  AOI21_X1  g754(.A(KEYINPUT126), .B1(new_n952_), .B2(new_n918_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n918_), .ZN(new_n957_));
  NOR4_X1   g756(.A1(new_n855_), .A2(new_n950_), .A3(new_n900_), .A4(new_n957_), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n692_), .B(new_n945_), .C1(new_n956_), .C2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n955_), .A2(new_n960_), .ZN(G1352gat));
  INV_X1    g760(.A(G204gat), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n954_), .A2(new_n962_), .A3(new_n651_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n651_), .B1(new_n956_), .B2(new_n958_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(G204gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n965_), .ZN(G1353gat));
  OR2_X1    g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n967_), .B1(new_n954_), .B2(new_n886_), .ZN(new_n968_));
  XOR2_X1   g767(.A(KEYINPUT63), .B(G211gat), .Z(new_n969_));
  OAI211_X1 g768(.A(new_n886_), .B(new_n969_), .C1(new_n956_), .C2(new_n958_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n968_), .A2(new_n971_), .ZN(G1354gat));
  NAND3_X1  g771(.A1(new_n954_), .A2(new_n360_), .A3(new_n253_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n257_), .B1(new_n951_), .B2(new_n953_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n360_), .B2(new_n974_), .ZN(G1355gat));
endmodule


