//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT72), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G85gat), .B(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(KEYINPUT64), .A3(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n212_), .A2(KEYINPUT65), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT65), .B1(new_n212_), .B2(new_n218_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT71), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n221_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n210_), .B(KEYINPUT69), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n232_), .B1(new_n224_), .B2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT8), .B1(new_n232_), .B2(KEYINPUT68), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT12), .B(new_n209_), .C1(new_n231_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n221_), .A2(new_n227_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n208_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT12), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n245_), .A2(new_n246_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G230gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n256_), .A3(new_n247_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n245_), .A2(KEYINPUT70), .A3(new_n246_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G120gat), .B(G148gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G176gat), .B(G204gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n262_), .B(new_n263_), .Z(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n255_), .A2(new_n259_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n255_), .B2(new_n259_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT13), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT75), .B(G43gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G50gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G29gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G15gat), .B(G22gat), .ZN(new_n276_));
  INV_X1    g075(.A(G1gat), .ZN(new_n277_));
  INV_X1    g076(.A(G8gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT14), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G8gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  AND2_X1   g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT15), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n275_), .B(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n284_), .B1(new_n286_), .B2(new_n282_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G229gat), .A2(G233gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n275_), .B(new_n282_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G113gat), .B(G141gat), .ZN(new_n293_));
  INV_X1    g092(.A(G169gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G197gat), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(KEYINPUT77), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n292_), .B(new_n297_), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n271_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT90), .ZN(new_n301_));
  INV_X1    g100(.A(G204gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT89), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT89), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G204gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(G197gat), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G197gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT21), .B1(new_n307_), .B2(new_n302_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n301_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT21), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(G204gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT89), .B(G204gat), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n311_), .B(new_n312_), .C1(new_n313_), .C2(new_n307_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(G197gat), .B2(G204gat), .ZN(new_n315_));
  OAI211_X1 g114(.A(KEYINPUT90), .B(new_n315_), .C1(new_n313_), .C2(G197gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n309_), .A2(new_n310_), .A3(new_n314_), .A4(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n310_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n311_), .B1(new_n318_), .B2(KEYINPUT91), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n310_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n312_), .B1(new_n313_), .B2(new_n307_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT22), .B(G169gat), .ZN(new_n326_));
  INV_X1    g125(.A(G176gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT23), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(G183gat), .A3(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n328_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n340_));
  NAND2_X1  g139(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n294_), .A2(new_n327_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n340_), .A2(new_n346_), .A3(new_n347_), .A4(new_n341_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n330_), .A2(new_n332_), .A3(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n331_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n336_), .B1(new_n345_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n324_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT22), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G169gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n294_), .A2(KEYINPUT22), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT79), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT79), .B1(new_n294_), .B2(KEYINPUT22), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n327_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n355_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(G176gat), .B1(new_n357_), .B2(KEYINPUT79), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n363_), .B(KEYINPUT80), .C1(KEYINPUT79), .C2(new_n326_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n350_), .A2(new_n351_), .A3(new_n334_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n347_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT24), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n343_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n333_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n325_), .A2(new_n343_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n337_), .A2(new_n338_), .B1(new_n372_), .B2(KEYINPUT24), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n333_), .A2(KEYINPUT78), .A3(new_n368_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n366_), .A2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n354_), .B(KEYINPUT20), .C1(new_n324_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT19), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT95), .B1(new_n324_), .B2(new_n353_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n353_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT95), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n323_), .A4(new_n317_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT20), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT94), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n376_), .A2(new_n324_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n376_), .B2(new_n324_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n380_), .B1(new_n387_), .B2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G8gat), .B(G36gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G64gat), .B(G92gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n376_), .A2(new_n324_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT94), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n389_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n405_), .A3(new_n386_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n380_), .A3(new_n398_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT27), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT101), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT101), .ZN(new_n412_));
  AOI211_X1 g211(.A(new_n412_), .B(KEYINPUT27), .C1(new_n400_), .C2(new_n407_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416_));
  INV_X1    g215(.A(G141gat), .ZN(new_n417_));
  INV_X1    g216(.A(G148gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n420_));
  NOR2_X1   g219(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G141gat), .A2(G148gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT2), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT2), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(G141gat), .A3(G148gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n422_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT88), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT88), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n422_), .A2(new_n427_), .A3(new_n432_), .A4(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G155gat), .ZN(new_n435_));
  INV_X1    g234(.A(G162gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G155gat), .A2(G162gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(G155gat), .B2(G162gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT86), .B1(new_n442_), .B2(new_n438_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444_));
  INV_X1    g243(.A(new_n438_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n444_), .B(new_n445_), .C1(new_n437_), .C2(new_n441_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n437_), .A2(new_n441_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n423_), .A3(new_n419_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n416_), .B1(new_n440_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n324_), .ZN(new_n451_));
  OAI211_X1 g250(.A(G228gat), .B(G233gat), .C1(new_n450_), .C2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n448_), .A2(new_n423_), .A3(new_n419_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n439_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n453_), .B(new_n324_), .C1(new_n457_), .C2(new_n416_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G78gat), .B(G106gat), .Z(new_n461_));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G22gat), .B(G50gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT28), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n440_), .A2(new_n449_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(KEYINPUT29), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(new_n416_), .A3(new_n464_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n462_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n460_), .A2(new_n461_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n461_), .B1(new_n452_), .B2(new_n458_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n472_), .B2(new_n469_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n460_), .A2(new_n461_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n471_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n377_), .A2(new_n379_), .ZN(new_n478_));
  OAI221_X1 g277(.A(KEYINPUT20), .B1(new_n324_), .B2(new_n353_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n379_), .ZN(new_n480_));
  OAI211_X1 g279(.A(KEYINPUT27), .B(new_n407_), .C1(new_n480_), .C2(new_n398_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n415_), .A2(KEYINPUT102), .A3(new_n477_), .A4(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n477_), .B(new_n481_), .C1(new_n410_), .C2(new_n413_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT102), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G15gat), .B(G43gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G71gat), .B(G99gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G227gat), .A2(G233gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT82), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n489_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n376_), .B(KEYINPUT30), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(KEYINPUT83), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n495_));
  OR2_X1    g294(.A1(G127gat), .A2(G134gat), .ZN(new_n496_));
  INV_X1    g295(.A(G113gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G127gat), .A2(G134gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G120gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n497_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n496_), .A2(new_n498_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G113gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(G120gat), .B1(new_n505_), .B2(new_n499_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n495_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n501_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(G120gat), .A3(new_n499_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(KEYINPUT84), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n494_), .B(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n493_), .A2(KEYINPUT83), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n512_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT0), .B(G57gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G85gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(G1gat), .B(G29gat), .Z(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n510_), .B(new_n507_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n503_), .A2(new_n506_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n440_), .A2(new_n523_), .A3(new_n449_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(KEYINPUT4), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G225gat), .A2(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT4), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n466_), .A2(new_n528_), .A3(new_n510_), .A4(new_n507_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n522_), .A2(new_n526_), .A3(new_n524_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n521_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n522_), .A2(KEYINPUT4), .A3(new_n524_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n527_), .B1(new_n522_), .B2(KEYINPUT4), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n531_), .B(new_n521_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n516_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n486_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n406_), .A2(new_n380_), .A3(new_n398_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n398_), .B1(new_n406_), .B2(new_n380_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n522_), .A2(new_n527_), .A3(new_n524_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n520_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n529_), .A2(new_n526_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n546_), .B2(new_n525_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(KEYINPUT33), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n536_), .A2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n530_), .A2(new_n531_), .A3(new_n521_), .A4(new_n549_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n547_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n400_), .A2(KEYINPUT97), .A3(new_n407_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n543_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n398_), .A2(KEYINPUT32), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n406_), .A2(new_n380_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n536_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n532_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n480_), .A2(new_n556_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT99), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n402_), .A2(new_n389_), .B1(new_n451_), .B2(new_n382_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n386_), .B1(new_n562_), .B2(KEYINPUT20), .ZN(new_n563_));
  OAI211_X1 g362(.A(KEYINPUT32), .B(new_n398_), .C1(new_n563_), .C2(new_n478_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT99), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n537_), .A2(new_n564_), .A3(new_n565_), .A4(new_n557_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n555_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n567_), .A2(KEYINPUT100), .A3(new_n477_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT100), .B1(new_n567_), .B2(new_n477_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n461_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n459_), .A2(new_n570_), .A3(new_n473_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n472_), .A2(new_n469_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n476_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n537_), .B1(new_n573_), .B2(new_n470_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n574_), .B(new_n481_), .C1(new_n410_), .C2(new_n413_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n568_), .A2(new_n569_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n516_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n539_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n300_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n282_), .B(new_n208_), .ZN(new_n581_));
  AND2_X1   g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT16), .B(G183gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT72), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT17), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(KEYINPUT17), .B2(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n583_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G134gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(new_n436_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT34), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n231_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n242_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n286_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n275_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n245_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n603_), .A2(new_n605_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n606_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NOR4_X1   g413(.A1(new_n609_), .A2(new_n603_), .A3(new_n605_), .A4(new_n611_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n600_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n231_), .A2(new_n242_), .ZN(new_n617_));
  OAI221_X1 g416(.A(new_n613_), .B1(new_n245_), .B2(new_n610_), .C1(new_n617_), .C2(new_n286_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n612_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n598_), .B(new_n599_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT37), .B1(new_n623_), .B2(KEYINPUT76), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT76), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT37), .ZN(new_n626_));
  AOI211_X1 g425(.A(new_n625_), .B(new_n626_), .C1(new_n616_), .C2(new_n622_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n580_), .A2(new_n595_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n277_), .A3(new_n537_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT38), .ZN(new_n631_));
  INV_X1    g430(.A(new_n580_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n623_), .B(KEYINPUT103), .Z(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(new_n594_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n537_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n631_), .A2(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(new_n481_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n634_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G8gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n629_), .A2(new_n278_), .A3(new_n641_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n645_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n642_), .A2(G8gat), .A3(new_n648_), .A4(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(KEYINPUT40), .A3(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n635_), .B2(new_n516_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT41), .Z(new_n660_));
  INV_X1    g459(.A(G15gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n629_), .A2(new_n661_), .A3(new_n578_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n635_), .B2(new_n477_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n477_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n629_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(G1327gat));
  NOR3_X1   g468(.A1(new_n580_), .A2(new_n633_), .A3(new_n594_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n537_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n579_), .A2(new_n672_), .A3(new_n628_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT106), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n567_), .A2(new_n477_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n567_), .A2(KEYINPUT100), .A3(new_n477_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n575_), .A3(new_n678_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n679_), .A2(new_n516_), .B1(new_n486_), .B2(new_n538_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n624_), .A2(new_n627_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n516_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n683_), .B2(new_n539_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n672_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n674_), .A2(new_n682_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT107), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n687_), .A2(new_n595_), .A3(new_n300_), .A4(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n688_), .A2(KEYINPUT107), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n690_), .A2(new_n691_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n636_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n671_), .B1(new_n695_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n670_), .A2(new_n697_), .A3(new_n641_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT108), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n670_), .A2(new_n700_), .A3(new_n697_), .A4(new_n641_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n699_), .A2(KEYINPUT45), .A3(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT45), .B1(new_n699_), .B2(new_n701_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n300_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n685_), .B1(new_n684_), .B2(new_n672_), .ZN(new_n706_));
  NOR4_X1   g505(.A1(new_n680_), .A2(KEYINPUT106), .A3(KEYINPUT43), .A4(new_n681_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n705_), .B1(new_n708_), .B2(new_n682_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n691_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n709_), .A2(new_n595_), .A3(new_n710_), .A4(new_n689_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n690_), .A2(new_n691_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n640_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n704_), .B1(new_n713_), .B2(new_n697_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n704_), .B(KEYINPUT46), .C1(new_n713_), .C2(new_n697_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n578_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G43gat), .ZN(new_n721_));
  INV_X1    g520(.A(G43gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n670_), .A2(new_n722_), .A3(new_n578_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n516_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n719_), .B(new_n723_), .C1(new_n725_), .C2(new_n722_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n724_), .A2(new_n727_), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n670_), .B2(new_n667_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n694_), .A2(new_n477_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G50gat), .ZN(G1331gat));
  NOR3_X1   g530(.A1(new_n680_), .A2(new_n299_), .A3(new_n271_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(new_n634_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n636_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n628_), .A2(new_n595_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n732_), .A2(new_n737_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT109), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT109), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n537_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n736_), .B1(new_n741_), .B2(new_n735_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n733_), .B2(new_n641_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT48), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n641_), .A2(new_n743_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n738_), .B2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n734_), .B2(new_n516_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n738_), .A2(G71gat), .A3(new_n516_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT110), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n733_), .B2(new_n667_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT50), .Z(new_n755_));
  NOR2_X1   g554(.A1(new_n477_), .A2(G78gat), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT111), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n738_), .B2(new_n757_), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n633_), .A2(new_n594_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n732_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n537_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n271_), .A2(new_n594_), .A3(new_n299_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n687_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n217_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n215_), .A2(new_n216_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n537_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT113), .Z(new_n769_));
  AOI21_X1  g568(.A(new_n763_), .B1(new_n765_), .B2(new_n769_), .ZN(G1336gat));
  AOI21_X1  g569(.A(G92gat), .B1(new_n762_), .B2(new_n641_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n765_), .A2(new_n641_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(G92gat), .B2(new_n772_), .ZN(G1337gat));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n226_), .A3(new_n578_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT114), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n765_), .A2(new_n578_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G99gat), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n762_), .A2(new_n778_), .A3(new_n226_), .A4(new_n578_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g580(.A1(new_n765_), .A2(new_n667_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT52), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(G106gat), .A3(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(KEYINPUT52), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n762_), .A2(new_n225_), .A3(new_n667_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n786_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n782_), .A2(G106gat), .A3(new_n789_), .A4(new_n784_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n787_), .A2(new_n793_), .A3(new_n788_), .A4(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n287_), .A2(new_n289_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n291_), .A2(new_n289_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n296_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n254_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n251_), .A2(new_n801_), .A3(new_n253_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n264_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT56), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n264_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n266_), .A3(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n800_), .B1(new_n809_), .B2(new_n298_), .ZN(new_n810_));
  OR2_X1    g609(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n810_), .A2(new_n633_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n810_), .B2(new_n633_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n806_), .A2(new_n266_), .A3(new_n799_), .A4(new_n808_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n628_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT119), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n815_), .A2(new_n816_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(new_n628_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n814_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n595_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n298_), .A2(new_n594_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n271_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n681_), .B1(new_n828_), .B2(new_n827_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OR3_X1    g632(.A1(new_n830_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n825_), .A2(new_n826_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n594_), .B1(new_n814_), .B2(new_n823_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT120), .B1(new_n839_), .B2(new_n836_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n486_), .A2(new_n537_), .A3(new_n578_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(KEYINPUT121), .Z(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n299_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n825_), .A2(new_n837_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n842_), .B(KEYINPUT123), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n846_), .A2(new_n299_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n845_), .B1(new_n851_), .B2(G113gat), .ZN(G1340gat));
  NAND2_X1  g651(.A1(new_n846_), .A2(new_n850_), .ZN(new_n853_));
  OAI21_X1  g652(.A(G120gat), .B1(new_n853_), .B2(new_n271_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n501_), .B1(new_n271_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n844_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n501_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1341gat));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT124), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n860_));
  OAI21_X1  g659(.A(G127gat), .B1(new_n595_), .B2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n846_), .A2(new_n850_), .A3(new_n859_), .A4(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n858_), .B1(new_n843_), .B2(new_n595_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n862_), .A2(KEYINPUT125), .A3(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1342gat));
  NOR2_X1   g667(.A1(new_n843_), .A2(new_n633_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(G134gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n853_), .A2(new_n681_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(G134gat), .ZN(G1343gat));
  AND2_X1   g671(.A1(new_n838_), .A2(new_n840_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n641_), .A2(new_n636_), .A3(new_n477_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n516_), .A3(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n298_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n417_), .ZN(G1344gat));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n271_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n418_), .ZN(G1345gat));
  NOR2_X1   g678(.A1(new_n875_), .A2(new_n595_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G155gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT126), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n880_), .B(new_n883_), .ZN(G1346gat));
  NOR3_X1   g683(.A1(new_n875_), .A2(new_n436_), .A3(new_n681_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n875_), .A2(new_n633_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n436_), .B2(new_n886_), .ZN(G1347gat));
  NAND2_X1  g686(.A1(new_n641_), .A2(new_n538_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n847_), .A2(new_n477_), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n298_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n294_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT62), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n326_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(KEYINPUT62), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(G1348gat));
  AND2_X1   g695(.A1(new_n873_), .A2(new_n477_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n271_), .A2(new_n327_), .A3(new_n888_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n890_), .A2(new_n271_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n897_), .A2(new_n898_), .B1(new_n899_), .B2(new_n327_), .ZN(G1349gat));
  NOR3_X1   g699(.A1(new_n890_), .A2(new_n595_), .A3(new_n337_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n897_), .A2(new_n594_), .A3(new_n889_), .ZN(new_n902_));
  INV_X1    g701(.A(G183gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n890_), .B2(new_n681_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n338_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n633_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n890_), .B2(new_n907_), .ZN(G1351gat));
  NOR3_X1   g707(.A1(new_n640_), .A2(new_n537_), .A3(new_n477_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n873_), .A2(new_n516_), .A3(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n298_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n307_), .ZN(G1352gat));
  OAI21_X1  g711(.A(G204gat), .B1(new_n910_), .B2(new_n271_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n910_), .A2(new_n271_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n313_), .ZN(G1353gat));
  NAND2_X1  g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n594_), .A2(new_n916_), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT127), .Z(new_n918_));
  NOR2_X1   g717(.A1(new_n910_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1354gat));
  INV_X1    g720(.A(G218gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n910_), .A2(new_n922_), .A3(new_n681_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n910_), .A2(new_n633_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(new_n924_), .ZN(G1355gat));
endmodule


