//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_, new_n999_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G43gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G50gat), .ZN(new_n206_));
  INV_X1    g005(.A(G43gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G50gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n206_), .A2(new_n210_), .A3(KEYINPUT15), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT15), .B1(new_n206_), .B2(new_n210_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  NOR2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n214_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT8), .B1(new_n214_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n221_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT64), .B(G106gat), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n227_), .A3(KEYINPUT65), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n214_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G85gat), .ZN(new_n236_));
  INV_X1    g035(.A(G92gat), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(KEYINPUT9), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n220_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n232_), .A2(new_n235_), .A3(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT67), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n239_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(new_n235_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n225_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT74), .B1(new_n213_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT34), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT35), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(KEYINPUT35), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n241_), .A2(KEYINPUT67), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n244_), .A2(new_n243_), .A3(new_n235_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n224_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n206_), .A2(new_n210_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .A4(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT15), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n208_), .A2(new_n209_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n205_), .A2(G50gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n206_), .A2(new_n210_), .A3(KEYINPUT15), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n258_), .B(new_n256_), .C1(new_n264_), .C2(new_n254_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT35), .A3(new_n249_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n257_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT75), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G190gat), .B(G218gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(G134gat), .ZN(new_n270_));
  INV_X1    g069(.A(G162gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT36), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT75), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n257_), .A2(new_n266_), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT36), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n267_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT37), .B1(new_n276_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT76), .B(G15gat), .ZN(new_n282_));
  INV_X1    g081(.A(G22gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G8gat), .ZN(new_n285_));
  INV_X1    g084(.A(G1gat), .ZN(new_n286_));
  INV_X1    g085(.A(G8gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT14), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n285_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n285_), .B1(new_n284_), .B2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT77), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(new_n289_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT78), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(new_n295_), .A3(KEYINPUT78), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G57gat), .B(G64gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G71gat), .B(G78gat), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n301_), .A2(KEYINPUT11), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n303_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n300_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G183gat), .B(G211gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G127gat), .B(G155gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n315_), .A2(KEYINPUT17), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n317_), .A3(KEYINPUT17), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n310_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n310_), .A2(new_n318_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT37), .ZN(new_n324_));
  INV_X1    g123(.A(new_n273_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n257_), .B2(new_n266_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n279_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n281_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n328_), .B(KEYINPUT80), .Z(new_n329_));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G78gat), .B(G106gat), .ZN(new_n331_));
  INV_X1    g130(.A(G155gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(new_n271_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G141gat), .ZN(new_n336_));
  INV_X1    g135(.A(G148gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT3), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(G141gat), .B2(G148gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT2), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n341_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n335_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT1), .B1(new_n332_), .B2(new_n271_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G155gat), .A3(G162gat), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n351_), .B(new_n353_), .C1(G155gat), .C2(G162gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n336_), .A2(new_n337_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n342_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n350_), .A2(KEYINPUT90), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT90), .B1(new_n350_), .B2(new_n356_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT29), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  INV_X1    g159(.A(G204gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT92), .ZN(new_n363_));
  INV_X1    g162(.A(G197gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(G204gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(G204gat), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n360_), .B(new_n362_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G211gat), .B(G218gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n361_), .A3(G197gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT91), .B1(new_n364_), .B2(G204gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n361_), .A2(G197gat), .ZN(new_n373_));
  OAI211_X1 g172(.A(KEYINPUT21), .B(new_n371_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n367_), .A2(new_n369_), .A3(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n362_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(KEYINPUT21), .A3(new_n368_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n359_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n350_), .B2(new_n356_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n378_), .ZN(new_n384_));
  OAI211_X1 g183(.A(G228gat), .B(G233gat), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n331_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n387_));
  INV_X1    g186(.A(new_n335_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n341_), .A2(new_n346_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT89), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n341_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n388_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n356_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n387_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n350_), .A2(KEYINPUT90), .A3(new_n356_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n382_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n380_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n385_), .B(new_n331_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n330_), .B1(new_n386_), .B2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n385_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n331_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(KEYINPUT93), .A3(new_n398_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n394_), .A2(new_n382_), .A3(new_n395_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G50gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT28), .B(G22gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n394_), .A2(new_n382_), .A3(new_n209_), .A4(new_n395_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n400_), .A2(new_n404_), .A3(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n386_), .A2(new_n399_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n406_), .A2(new_n409_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n407_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n410_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n418_), .A3(KEYINPUT93), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n421_));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n427_));
  NAND2_X1  g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428_));
  INV_X1    g227(.A(G169gat), .ZN(new_n429_));
  INV_X1    g228(.A(G176gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n428_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G183gat), .A2(G190gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT23), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT23), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G183gat), .A3(G190gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT26), .B(G190gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT25), .B(G183gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n432_), .A2(new_n437_), .A3(new_n440_), .A4(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(G183gat), .ZN(new_n444_));
  INV_X1    g243(.A(G190gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n437_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT22), .B(G169gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n430_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n428_), .B(KEYINPUT95), .ZN(new_n450_));
  AND4_X1   g249(.A1(KEYINPUT96), .A2(new_n447_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n437_), .A2(new_n446_), .B1(new_n448_), .B2(new_n430_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT96), .B1(new_n452_), .B2(new_n450_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n443_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n378_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n456_));
  NOR3_X1   g255(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n457_), .B(new_n459_), .C1(new_n437_), .C2(new_n446_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT84), .B(KEYINPUT26), .C1(new_n445_), .C2(KEYINPUT85), .ZN(new_n461_));
  NAND2_X1  g260(.A1(KEYINPUT84), .A2(KEYINPUT26), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(G190gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT26), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(G190gat), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n461_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n444_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n444_), .B2(KEYINPUT83), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n470_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n469_), .B(KEYINPUT25), .C1(new_n444_), .C2(KEYINPUT83), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n468_), .A2(new_n472_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n431_), .A2(KEYINPUT24), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n431_), .A2(KEYINPUT24), .A3(new_n428_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n437_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n460_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n456_), .B1(new_n481_), .B2(new_n384_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT19), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n455_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n474_), .A2(new_n475_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n461_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n471_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n447_), .A2(new_n458_), .ZN(new_n489_));
  OAI22_X1  g288(.A1(new_n488_), .A2(new_n479_), .B1(new_n457_), .B2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n456_), .B1(new_n490_), .B2(new_n378_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n384_), .B(new_n443_), .C1(new_n453_), .C2(new_n451_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n484_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n426_), .B1(new_n485_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n484_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n454_), .A2(new_n378_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT20), .B1(new_n481_), .B2(new_n384_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n455_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n425_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n494_), .A2(KEYINPUT98), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT27), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT98), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n503_), .B(new_n426_), .C1(new_n485_), .C2(new_n493_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n452_), .A2(new_n450_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n443_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n508_), .B2(new_n378_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT102), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n509_), .A2(KEYINPUT102), .B1(new_n378_), .B2(new_n490_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n495_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n455_), .A2(new_n482_), .A3(new_n495_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(KEYINPUT27), .B(new_n494_), .C1(new_n514_), .C2(new_n426_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n505_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n420_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G120gat), .ZN(new_n519_));
  AND2_X1   g318(.A1(G127gat), .A2(G134gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G127gat), .A2(G134gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT87), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(G127gat), .ZN(new_n523_));
  INV_X1    g322(.A(G134gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G127gat), .A2(G134gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(G113gat), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n522_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n529_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n519_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n522_), .A2(new_n528_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(G113gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n522_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(G120gat), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G225gat), .A2(G233gat), .ZN(new_n539_));
  AND4_X1   g338(.A1(new_n350_), .A2(new_n532_), .A3(new_n536_), .A4(new_n356_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT100), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n394_), .A2(new_n395_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n540_), .B1(new_n545_), .B2(new_n537_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(KEYINPUT100), .A3(new_n539_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n549_));
  XNOR2_X1  g348(.A(G1gat), .B(G29gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G57gat), .B(G85gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n539_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT4), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n532_), .A2(new_n536_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(KEYINPUT4), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n554_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n548_), .A2(new_n553_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n553_), .B1(new_n548_), .B2(new_n560_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT86), .B(G99gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G43gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n537_), .B(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G227gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n481_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT30), .B(G71gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n569_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n563_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n518_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n505_), .A2(new_n515_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n420_), .A2(KEYINPUT104), .A3(new_n578_), .A4(new_n563_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT104), .ZN(new_n580_));
  INV_X1    g379(.A(new_n553_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT100), .B1(new_n546_), .B2(new_n539_), .ZN(new_n582_));
  NOR4_X1   g381(.A1(new_n558_), .A2(new_n543_), .A3(new_n554_), .A4(new_n540_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT4), .B1(new_n558_), .B2(new_n540_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n538_), .A2(new_n555_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n539_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n581_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n548_), .A2(new_n553_), .A3(new_n560_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n414_), .A2(new_n588_), .A3(new_n419_), .A4(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n580_), .B1(new_n590_), .B2(new_n516_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n579_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n512_), .A2(new_n513_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(new_n593_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT103), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n588_), .A2(new_n589_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT103), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n596_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n589_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n501_), .A2(new_n504_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n539_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n546_), .A2(new_n554_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n581_), .A3(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n548_), .A2(new_n560_), .A3(KEYINPUT33), .A4(new_n553_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n603_), .A2(new_n604_), .A3(new_n607_), .A4(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n598_), .A2(new_n601_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n420_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n592_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n577_), .B1(new_n613_), .B2(new_n574_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n255_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n298_), .A2(new_n617_), .A3(new_n299_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n299_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT78), .B1(new_n292_), .B2(new_n295_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n213_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n300_), .A2(new_n255_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n615_), .A3(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G113gat), .B(G141gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT81), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(G169gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(new_n364_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n621_), .A2(new_n627_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n627_), .B2(new_n621_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n307_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n246_), .A2(KEYINPUT69), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n636_), .A2(KEYINPUT69), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(KEYINPUT69), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n254_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n637_), .A2(new_n639_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT70), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT12), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(KEYINPUT71), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n246_), .A2(new_n646_), .A3(new_n307_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n646_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n636_), .B1(new_n254_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n254_), .A2(new_n645_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n647_), .A2(new_n649_), .A3(new_n638_), .A4(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT70), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n637_), .A2(new_n642_), .A3(new_n652_), .A4(new_n639_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n644_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n657_), .B(new_n658_), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n654_), .B(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT13), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n614_), .A2(new_n635_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n329_), .A2(new_n666_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n667_), .A2(G1gat), .A3(new_n563_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n579_), .A2(new_n591_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n611_), .B2(new_n610_), .ZN(new_n675_));
  OAI22_X1  g474(.A1(new_n675_), .A2(new_n575_), .B1(new_n518_), .B2(new_n576_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n257_), .A2(new_n266_), .A3(new_n274_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n274_), .B1(new_n257_), .B2(new_n266_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n325_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n279_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(KEYINPUT106), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(new_n614_), .B2(new_n680_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n682_), .A2(new_n684_), .A3(new_n322_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n665_), .A2(new_n635_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G1gat), .B1(new_n687_), .B2(new_n563_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n672_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n673_), .A2(new_n688_), .A3(new_n689_), .ZN(G1324gat));
  INV_X1    g489(.A(new_n667_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n287_), .A3(new_n516_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n685_), .A2(new_n686_), .A3(new_n516_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT39), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(G8gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n693_), .B2(G8gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n692_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT40), .B(new_n692_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1325gat));
  OR3_X1    g501(.A1(new_n667_), .A2(G15gat), .A3(new_n574_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n685_), .A2(new_n686_), .A3(new_n575_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT41), .B1(new_n704_), .B2(G15gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(G1326gat));
  NAND3_X1  g507(.A1(new_n691_), .A2(new_n283_), .A3(new_n420_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n685_), .A2(new_n686_), .A3(new_n420_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(G22gat), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n710_), .B2(G22gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n713_), .B2(new_n714_), .ZN(G1327gat));
  NOR2_X1   g514(.A1(new_n681_), .A2(new_n322_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n666_), .A2(new_n716_), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n717_), .A2(G29gat), .A3(new_n563_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n686_), .A2(new_n323_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n324_), .B1(new_n679_), .B2(new_n279_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n327_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n676_), .B2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n575_), .B1(new_n592_), .B2(new_n612_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n721_), .B(new_n724_), .C1(new_n726_), .C2(new_n577_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n720_), .B1(new_n725_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n724_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n614_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n719_), .B1(new_n733_), .B2(new_n727_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT44), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n599_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT107), .B1(new_n736_), .B2(G29gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n599_), .B1(new_n734_), .B2(KEYINPUT44), .ZN(new_n738_));
  AOI211_X1 g537(.A(new_n730_), .B(new_n719_), .C1(new_n733_), .C2(new_n727_), .ZN(new_n739_));
  OAI211_X1 g538(.A(KEYINPUT107), .B(G29gat), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n718_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT108), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n718_), .C1(new_n737_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1328gat));
  INV_X1    g545(.A(G36gat), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n676_), .A2(new_n686_), .A3(new_n747_), .A4(new_n716_), .ZN(new_n748_));
  OR3_X1    g547(.A1(new_n748_), .A2(KEYINPUT109), .A3(new_n578_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT109), .B1(new_n748_), .B2(new_n578_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n739_), .A2(new_n578_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n747_), .B1(new_n755_), .B2(new_n731_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n758_));
  OR2_X1    g557(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n754_), .A2(new_n757_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n752_), .A2(new_n753_), .ZN(new_n761_));
  OAI211_X1 g560(.A(KEYINPUT110), .B(KEYINPUT46), .C1(new_n761_), .C2(new_n756_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1329gat));
  OAI21_X1  g562(.A(new_n207_), .B1(new_n717_), .B2(new_n574_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n735_), .A2(G43gat), .A3(new_n575_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n731_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g567(.A(new_n717_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G50gat), .B1(new_n769_), .B2(new_n420_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n766_), .A2(new_n739_), .A3(new_n209_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n420_), .ZN(G1331gat));
  INV_X1    g571(.A(G57gat), .ZN(new_n773_));
  INV_X1    g572(.A(new_n635_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n663_), .A2(new_n664_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n614_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n329_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n777_), .B2(new_n563_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT111), .Z(new_n779_));
  NOR2_X1   g578(.A1(new_n775_), .A2(new_n774_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n685_), .A2(G57gat), .A3(new_n599_), .A4(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1332gat));
  OR3_X1    g581(.A1(new_n777_), .A2(G64gat), .A3(new_n578_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n685_), .A2(new_n516_), .A3(new_n780_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT48), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(G64gat), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n784_), .B2(G64gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n783_), .B1(new_n787_), .B2(new_n788_), .ZN(G1333gat));
  OR3_X1    g588(.A1(new_n777_), .A2(G71gat), .A3(new_n574_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n685_), .A2(new_n575_), .A3(new_n780_), .ZN(new_n791_));
  XOR2_X1   g590(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(G71gat), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n791_), .B2(G71gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n790_), .B1(new_n794_), .B2(new_n795_), .ZN(G1334gat));
  OR3_X1    g595(.A1(new_n777_), .A2(G78gat), .A3(new_n611_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n685_), .A2(new_n420_), .A3(new_n780_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(G78gat), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n798_), .B2(G78gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n797_), .B1(new_n801_), .B2(new_n802_), .ZN(G1335gat));
  NAND2_X1  g602(.A1(new_n776_), .A2(new_n716_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(G85gat), .B1(new_n805_), .B2(new_n599_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n780_), .A2(new_n323_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n733_), .B2(new_n727_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n563_), .A2(new_n236_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT113), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n806_), .B1(new_n808_), .B2(new_n810_), .ZN(G1336gat));
  AOI21_X1  g610(.A(G92gat), .B1(new_n805_), .B2(new_n516_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n578_), .A2(new_n237_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n808_), .B2(new_n813_), .ZN(G1337gat));
  INV_X1    g613(.A(new_n226_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n804_), .A2(new_n815_), .A3(new_n574_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT114), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n808_), .A2(new_n575_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G99gat), .ZN(new_n819_));
  AOI211_X1 g618(.A(KEYINPUT115), .B(KEYINPUT51), .C1(new_n817_), .C2(new_n819_), .ZN(new_n820_));
  OR2_X1    g619(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n821_));
  NAND2_X1  g620(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n822_));
  AND4_X1   g621(.A1(new_n821_), .A2(new_n817_), .A3(new_n822_), .A4(new_n819_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1338gat));
  NAND2_X1  g623(.A1(new_n808_), .A2(new_n420_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G106gat), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT116), .A3(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n805_), .A2(new_n227_), .A3(new_n420_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n827_), .A2(KEYINPUT116), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(KEYINPUT116), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n825_), .A2(G106gat), .A3(new_n830_), .A4(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n829_), .A3(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g633(.A1(new_n722_), .A2(new_n635_), .A3(new_n322_), .A4(new_n723_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT117), .B1(new_n835_), .B2(new_n665_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n328_), .A2(new_n837_), .A3(new_n635_), .A4(new_n775_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n838_), .A3(KEYINPUT54), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT117), .B(new_n840_), .C1(new_n835_), .C2(new_n665_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n654_), .A2(new_n660_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n647_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n639_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT55), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n651_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n844_), .A2(new_n848_), .A3(new_n639_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n659_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n843_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n616_), .B1(new_n626_), .B2(new_n618_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n632_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n615_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT119), .B1(new_n857_), .B2(new_n631_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n625_), .A2(new_n616_), .A3(new_n626_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n633_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n651_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(KEYINPUT55), .B2(new_n845_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n660_), .B1(new_n863_), .B2(new_n849_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT56), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n853_), .A2(new_n861_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n853_), .A2(new_n861_), .A3(KEYINPUT58), .A4(new_n865_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n724_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n852_), .B1(new_n851_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n843_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n864_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n872_), .A2(new_n774_), .A3(new_n873_), .A4(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n861_), .A2(new_n661_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n680_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n870_), .B1(KEYINPUT57), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n847_), .A2(new_n850_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n871_), .B1(new_n879_), .B2(new_n660_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n635_), .B1(new_n880_), .B2(KEYINPUT56), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n864_), .A2(KEYINPUT118), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n843_), .B1(new_n882_), .B2(new_n852_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n881_), .A2(new_n883_), .B1(new_n661_), .B2(new_n861_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885_));
  NOR4_X1   g684(.A1(new_n884_), .A2(KEYINPUT120), .A3(new_n885_), .A4(new_n680_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n877_), .B2(KEYINPUT57), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n878_), .A2(new_n886_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n842_), .B1(new_n889_), .B2(new_n322_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n563_), .A2(new_n574_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n517_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT59), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n890_), .A2(new_n894_), .A3(new_n517_), .A4(new_n891_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n893_), .A2(G113gat), .A3(new_n774_), .A4(new_n895_), .ZN(new_n896_));
  AND4_X1   g695(.A1(new_n774_), .A2(new_n890_), .A3(new_n517_), .A4(new_n891_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT121), .B1(new_n897_), .B2(G113gat), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n899_), .B(new_n529_), .C1(new_n892_), .C2(new_n635_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n896_), .A2(new_n898_), .A3(new_n900_), .ZN(G1340gat));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n775_), .B2(G120gat), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n890_), .A2(new_n517_), .A3(new_n891_), .A4(new_n903_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n893_), .A2(new_n665_), .A3(new_n895_), .A4(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G120gat), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n904_), .A2(KEYINPUT60), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1341gat));
  INV_X1    g707(.A(new_n892_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G127gat), .B1(new_n909_), .B2(new_n322_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n893_), .A2(new_n895_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n323_), .A2(new_n523_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1342gat));
  AOI21_X1  g712(.A(G134gat), .B1(new_n909_), .B2(new_n680_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n732_), .A2(new_n524_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n911_), .B2(new_n915_), .ZN(G1343gat));
  NAND2_X1  g715(.A1(new_n839_), .A2(new_n841_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n877_), .A2(KEYINPUT57), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT120), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n885_), .B1(new_n884_), .B2(new_n680_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n877_), .A2(new_n887_), .A3(KEYINPUT57), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n870_), .A4(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n917_), .B1(new_n922_), .B2(new_n323_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n611_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n563_), .A2(new_n575_), .A3(new_n516_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n924_), .A2(new_n774_), .A3(new_n925_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT122), .B(G141gat), .Z(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1344gat));
  AND2_X1   g727(.A1(new_n924_), .A2(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n665_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(G148gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n337_), .A3(new_n665_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1345gat));
  NAND3_X1  g732(.A1(new_n924_), .A2(new_n322_), .A3(new_n925_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT61), .B(G155gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1346gat));
  NAND2_X1  g735(.A1(new_n929_), .A2(new_n680_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n732_), .A2(new_n271_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n937_), .A2(new_n271_), .B1(new_n929_), .B2(new_n938_), .ZN(G1347gat));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n576_), .A2(new_n420_), .A3(new_n578_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n923_), .A2(new_n635_), .A3(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n940_), .B1(new_n943_), .B2(new_n429_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n890_), .A2(new_n774_), .A3(new_n941_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n945_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n944_), .A2(KEYINPUT62), .A3(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n943_), .A2(new_n448_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n940_), .B(new_n949_), .C1(new_n943_), .C2(new_n429_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n947_), .A2(new_n948_), .A3(new_n950_), .ZN(G1348gat));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n952_), .A2(G176gat), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n923_), .A2(new_n942_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n665_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n952_), .A2(G176gat), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n953_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n957_), .B1(new_n955_), .B2(new_n953_), .ZN(G1349gat));
  NAND2_X1  g757(.A1(new_n954_), .A2(new_n322_), .ZN(new_n959_));
  MUX2_X1   g758(.A(new_n439_), .B(G183gat), .S(new_n959_), .Z(G1350gat));
  NAND2_X1  g759(.A1(new_n680_), .A2(new_n438_), .ZN(new_n961_));
  XOR2_X1   g760(.A(new_n961_), .B(KEYINPUT125), .Z(new_n962_));
  NAND2_X1  g761(.A1(new_n954_), .A2(new_n962_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n923_), .A2(new_n732_), .A3(new_n942_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n964_), .B2(new_n445_), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  OAI211_X1 g766(.A(new_n963_), .B(KEYINPUT126), .C1(new_n445_), .C2(new_n964_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(G1351gat));
  INV_X1    g768(.A(new_n590_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n578_), .A2(new_n575_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n886_), .A2(new_n888_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n878_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n322_), .B1(new_n972_), .B2(new_n973_), .ZN(new_n974_));
  OAI211_X1 g773(.A(new_n970_), .B(new_n971_), .C1(new_n974_), .C2(new_n917_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  NAND4_X1  g776(.A1(new_n890_), .A2(KEYINPUT127), .A3(new_n970_), .A4(new_n971_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n977_), .A2(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(G197gat), .B1(new_n979_), .B2(new_n774_), .ZN(new_n980_));
  AOI211_X1 g779(.A(new_n364_), .B(new_n635_), .C1(new_n977_), .C2(new_n978_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n980_), .A2(new_n981_), .ZN(G1352gat));
  NAND2_X1  g781(.A1(new_n922_), .A2(new_n323_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n590_), .B1(new_n983_), .B2(new_n842_), .ZN(new_n984_));
  AOI21_X1  g783(.A(KEYINPUT127), .B1(new_n984_), .B2(new_n971_), .ZN(new_n985_));
  INV_X1    g784(.A(new_n971_), .ZN(new_n986_));
  NOR4_X1   g785(.A1(new_n923_), .A2(new_n976_), .A3(new_n590_), .A4(new_n986_), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n665_), .B1(new_n985_), .B2(new_n987_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n988_), .A2(G204gat), .ZN(new_n989_));
  NAND3_X1  g788(.A1(new_n979_), .A2(new_n361_), .A3(new_n665_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n989_), .A2(new_n990_), .ZN(G1353gat));
  OR2_X1    g790(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n992_));
  AOI21_X1  g791(.A(new_n992_), .B1(new_n979_), .B2(new_n322_), .ZN(new_n993_));
  XNOR2_X1  g792(.A(KEYINPUT63), .B(G211gat), .ZN(new_n994_));
  AOI211_X1 g793(.A(new_n323_), .B(new_n994_), .C1(new_n977_), .C2(new_n978_), .ZN(new_n995_));
  NOR2_X1   g794(.A1(new_n993_), .A2(new_n995_), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n979_), .B2(new_n680_), .ZN(new_n997_));
  INV_X1    g796(.A(G218gat), .ZN(new_n998_));
  AOI211_X1 g797(.A(new_n998_), .B(new_n732_), .C1(new_n977_), .C2(new_n978_), .ZN(new_n999_));
  NOR2_X1   g798(.A1(new_n997_), .A2(new_n999_), .ZN(G1355gat));
endmodule


