//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT93), .Z(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G197gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT92), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(new_n207_), .B2(new_n206_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(KEYINPUT21), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n202_), .B(KEYINPUT93), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT21), .B1(new_n206_), .B2(new_n205_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n211_), .B(new_n212_), .C1(new_n209_), .C2(KEYINPUT21), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G228gat), .A2(G233gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT87), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT2), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n219_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(new_n217_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229_));
  AND2_X1   g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G155gat), .ZN(new_n233_));
  INV_X1    g032(.A(G162gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT88), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n232_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT89), .B1(new_n228_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G141gat), .ZN(new_n240_));
  INV_X1    g039(.A(G148gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT87), .B1(new_n242_), .B2(KEYINPUT3), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n222_), .A2(KEYINPUT2), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n220_), .A2(G141gat), .A3(G148gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n243_), .A2(new_n246_), .A3(new_n225_), .A4(new_n219_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n232_), .A2(new_n237_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n242_), .A2(KEYINPUT85), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT85), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n216_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n222_), .A3(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n236_), .A2(KEYINPUT1), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n236_), .B1(new_n231_), .B2(KEYINPUT1), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT86), .B(new_n236_), .C1(new_n231_), .C2(KEYINPUT1), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n255_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n251_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT91), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT29), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n263_), .B2(KEYINPUT29), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n214_), .B(new_n215_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G78gat), .B(G106gat), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n215_), .B1(new_n272_), .B2(new_n214_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n268_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n214_), .A2(new_n215_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n263_), .A2(KEYINPUT29), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT91), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n278_), .B2(new_n265_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n269_), .B1(new_n279_), .B2(new_n273_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n263_), .B2(KEYINPUT29), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G22gat), .B(G50gat), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n261_), .B1(new_n239_), .B2(new_n250_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT29), .ZN(new_n285_));
  INV_X1    g084(.A(new_n281_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n282_), .A2(new_n283_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n282_), .B2(new_n287_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n275_), .A2(new_n280_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n275_), .B2(new_n280_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G8gat), .B(G36gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT18), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT20), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT26), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(G190gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(G190gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(KEYINPUT82), .B2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n302_), .A2(KEYINPUT82), .ZN(new_n304_));
  INV_X1    g103(.A(G183gat), .ZN(new_n305_));
  OR3_X1    g104(.A1(new_n305_), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT25), .B1(new_n305_), .B2(KEYINPUT81), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n303_), .A2(new_n304_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n309_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G183gat), .A3(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n321_), .B(new_n322_), .C1(G183gat), .C2(G190gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G169gat), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n308_), .A2(new_n319_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n299_), .B1(new_n214_), .B2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n210_), .A2(new_n213_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n318_), .B1(G183gat), .B2(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT95), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT95), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n333_), .A3(new_n325_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n321_), .A2(new_n322_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n301_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n302_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n338_), .A2(new_n313_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n332_), .A2(new_n334_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT19), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n328_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n332_), .A2(new_n334_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n339_), .A2(new_n335_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n299_), .B1(new_n349_), .B2(new_n214_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n326_), .A2(new_n213_), .A3(new_n210_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n344_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n298_), .B1(new_n346_), .B2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n351_), .B(KEYINPUT20), .C1(new_n329_), .C2(new_n340_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n343_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(new_n297_), .A3(new_n345_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n354_), .A2(new_n343_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n210_), .A2(new_n213_), .A3(new_n348_), .A4(new_n331_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n344_), .B1(new_n328_), .B2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n297_), .B(KEYINPUT101), .Z(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT27), .B(new_n356_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n359_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n293_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G127gat), .B(G134gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n369_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n368_), .A2(new_n369_), .A3(KEYINPUT84), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n284_), .A2(KEYINPUT4), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT96), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n370_), .A2(new_n372_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n284_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n249_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n262_), .B(new_n378_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT96), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n375_), .B1(new_n251_), .B2(new_n262_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n379_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n376_), .B1(new_n385_), .B2(KEYINPUT4), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n382_), .B(KEYINPUT96), .C1(new_n284_), .C2(new_n375_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n390_), .B2(new_n379_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G57gat), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n389_), .A2(new_n398_), .A3(new_n392_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403_));
  INV_X1    g202(.A(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n326_), .B(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(new_n375_), .Z(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(G15gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT30), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT31), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n407_), .B(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n402_), .A2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n367_), .A2(new_n414_), .ZN(new_n415_));
  AOI211_X1 g214(.A(new_n399_), .B(new_n391_), .C1(new_n386_), .C2(new_n388_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT33), .B1(new_n416_), .B2(KEYINPUT98), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT99), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n390_), .B2(new_n379_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n420_), .A2(new_n388_), .A3(new_n376_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n382_), .A2(KEYINPUT96), .ZN(new_n422_));
  INV_X1    g221(.A(new_n384_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n377_), .B1(new_n284_), .B2(new_n378_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n399_), .B1(new_n425_), .B2(new_n387_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n418_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n376_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n428_), .B(new_n387_), .C1(new_n425_), .C2(new_n419_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n398_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(KEYINPUT99), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n357_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n401_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n417_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT100), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n417_), .A2(new_n432_), .A3(KEYINPUT100), .A4(new_n435_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n270_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n279_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n440_), .A2(new_n441_), .B1(new_n289_), .B2(new_n288_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n275_), .A2(new_n280_), .A3(new_n290_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n355_), .A2(new_n345_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n297_), .A2(KEYINPUT32), .ZN(new_n446_));
  MUX2_X1   g245(.A(new_n363_), .B(new_n445_), .S(new_n446_), .Z(new_n447_));
  AOI21_X1  g246(.A(new_n398_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(new_n416_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n438_), .A2(new_n439_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n413_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n402_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n366_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n455_), .B2(new_n293_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n415_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n458_));
  XOR2_X1   g257(.A(G29gat), .B(G36gat), .Z(new_n459_));
  XOR2_X1   g258(.A(G43gat), .B(G50gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G1gat), .B(G8gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT76), .B(G15gat), .ZN(new_n464_));
  INV_X1    g263(.A(G22gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT77), .B(G8gat), .ZN(new_n467_));
  INV_X1    g266(.A(G1gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT14), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n463_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n469_), .A3(new_n463_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n462_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n472_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n474_), .A2(new_n461_), .A3(new_n470_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n458_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G229gat), .A2(G233gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n461_), .B1(new_n474_), .B2(new_n470_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(new_n462_), .A3(new_n472_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(KEYINPUT78), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(new_n478_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n462_), .A2(KEYINPUT15), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n461_), .A2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n483_), .A2(new_n471_), .A3(new_n485_), .A4(new_n472_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n477_), .B(KEYINPUT79), .Z(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(KEYINPUT80), .A3(new_n479_), .A4(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n479_), .A3(new_n487_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT80), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n482_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G169gat), .B(G197gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n482_), .A2(new_n488_), .A3(new_n491_), .A4(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n457_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G120gat), .B(G148gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT5), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G176gat), .B(G204gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G85gat), .B(G92gat), .ZN(new_n507_));
  INV_X1    g306(.A(G92gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(KEYINPUT9), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT65), .B(G85gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(new_n508_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT10), .B(G99gat), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT6), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT66), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT66), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT6), .ZN(new_n518_));
  AND2_X1   g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n521_));
  OAI221_X1 g320(.A(new_n513_), .B1(G106gat), .B2(new_n514_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT8), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT69), .B1(new_n520_), .B2(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n517_), .A2(KEYINPUT6), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n515_), .A2(KEYINPUT66), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT69), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(G99gat), .B2(G106gat), .ZN(new_n533_));
  INV_X1    g332(.A(G99gat), .ZN(new_n534_));
  INV_X1    g333(.A(G106gat), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n534_), .B(new_n535_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n524_), .A2(new_n531_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n507_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n523_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n523_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n537_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT68), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n537_), .B(new_n544_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n541_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n522_), .B1(new_n540_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G78gat), .Z(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n547_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT71), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n522_), .B(new_n554_), .C1(new_n540_), .C2(new_n546_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT70), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n547_), .A2(new_n560_), .A3(new_n555_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(KEYINPUT70), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n557_), .A2(new_n559_), .A3(new_n561_), .A4(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G230gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n556_), .A2(KEYINPUT12), .A3(new_n558_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n547_), .A2(new_n568_), .A3(new_n555_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n564_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n506_), .B1(new_n566_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n571_), .A3(new_n506_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(KEYINPUT13), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT13), .B1(new_n573_), .B2(new_n574_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n522_), .B(new_n461_), .C1(new_n540_), .C2(new_n546_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT35), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n483_), .A2(new_n485_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n547_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n583_), .A2(new_n584_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n586_), .B(new_n588_), .C1(KEYINPUT73), .C2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n579_), .A2(KEYINPUT73), .A3(new_n585_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n547_), .A2(new_n587_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n579_), .A2(new_n585_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n592_), .B(new_n589_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT36), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n591_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n598_), .B(KEYINPUT36), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT37), .B1(new_n601_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT74), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT74), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n607_), .B(KEYINPUT37), .C1(new_n601_), .C2(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n591_), .A2(new_n595_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n602_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n600_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n604_), .A2(new_n611_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n613_), .A2(KEYINPUT37), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n554_), .B(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n474_), .A2(new_n470_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G127gat), .B(G155gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT16), .ZN(new_n622_));
  XOR2_X1   g421(.A(G183gat), .B(G211gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT17), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n625_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n620_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n627_), .B2(new_n620_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n578_), .A2(new_n616_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n501_), .A2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(G1gat), .A3(new_n453_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(KEYINPUT104), .B2(KEYINPUT38), .ZN(new_n634_));
  NOR2_X1   g433(.A1(KEYINPUT104), .A2(KEYINPUT38), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n610_), .A2(new_n602_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT75), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n640_), .A2(KEYINPUT102), .A3(new_n600_), .A4(new_n612_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n457_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT103), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n578_), .A2(new_n630_), .A3(new_n500_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(new_n402_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n636_), .B1(new_n468_), .B2(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(new_n632_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n366_), .A3(new_n467_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(new_n366_), .A3(new_n645_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  AND4_X1   g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .A4(G8gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(G8gat), .B1(new_n651_), .B2(new_n653_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n652_), .A2(new_n656_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n650_), .B1(new_n654_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(G1325gat));
  AOI21_X1  g459(.A(new_n409_), .B1(new_n646_), .B2(new_n452_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT41), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n649_), .A2(new_n409_), .A3(new_n452_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  AOI21_X1  g463(.A(new_n465_), .B1(new_n646_), .B2(new_n293_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT42), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n649_), .A2(new_n465_), .A3(new_n293_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1327gat));
  NAND2_X1  g467(.A1(new_n642_), .A2(new_n630_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n578_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n501_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n402_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n609_), .A2(new_n615_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n457_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n402_), .A2(new_n366_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n413_), .B1(new_n676_), .B2(new_n444_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n444_), .A2(new_n449_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n437_), .B2(new_n436_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n679_), .B2(new_n439_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n675_), .B(new_n616_), .C1(new_n680_), .C2(new_n415_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n674_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n577_), .A2(new_n630_), .A3(new_n499_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n683_), .B1(new_n674_), .B2(new_n681_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n451_), .A2(new_n456_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n415_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n675_), .B1(new_n693_), .B2(new_n616_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n457_), .A2(KEYINPUT43), .A3(new_n673_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n684_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n687_), .A2(new_n689_), .B1(new_n690_), .B2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n402_), .A2(G29gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n672_), .B1(new_n697_), .B2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(G36gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n671_), .A2(new_n700_), .A3(new_n366_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT45), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n366_), .B1(new_n688_), .B2(KEYINPUT44), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n704_), .A2(KEYINPUT107), .A3(new_n700_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n454_), .B1(new_n696_), .B2(new_n690_), .ZN(new_n707_));
  AND4_X1   g506(.A1(KEYINPUT106), .A2(new_n682_), .A3(KEYINPUT44), .A4(new_n684_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT106), .B1(new_n688_), .B2(KEYINPUT44), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n706_), .B1(new_n710_), .B2(G36gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n702_), .B1(new_n705_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT46), .B(new_n702_), .C1(new_n705_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  NAND3_X1  g515(.A1(new_n697_), .A2(G43gat), .A3(new_n452_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n671_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n404_), .B1(new_n718_), .B2(new_n413_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g520(.A(G50gat), .B1(new_n671_), .B2(new_n293_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n293_), .A2(G50gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n697_), .B2(new_n723_), .ZN(G1331gat));
  INV_X1    g523(.A(G57gat), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n457_), .A2(new_n499_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n630_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n578_), .A4(new_n673_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n728_), .B2(new_n453_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT108), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n577_), .A2(new_n630_), .A3(new_n499_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n644_), .A2(new_n731_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n732_), .A2(KEYINPUT109), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(KEYINPUT109), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n453_), .A2(new_n725_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n730_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n366_), .A3(new_n734_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G64gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n454_), .A2(G64gat), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT110), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n740_), .A2(new_n741_), .B1(new_n728_), .B2(new_n743_), .ZN(G1333gat));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n452_), .A3(new_n734_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G71gat), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n413_), .A2(G71gat), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT111), .Z(new_n750_));
  OAI22_X1  g549(.A1(new_n747_), .A2(new_n748_), .B1(new_n728_), .B2(new_n750_), .ZN(G1334gat));
  OR3_X1    g550(.A1(new_n728_), .A2(G78gat), .A3(new_n444_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n733_), .A2(new_n293_), .A3(new_n734_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(G78gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G78gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1335gat));
  NOR2_X1   g556(.A1(new_n669_), .A2(new_n577_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n726_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n402_), .ZN(new_n761_));
  AND4_X1   g560(.A1(new_n630_), .A2(new_n682_), .A3(new_n500_), .A4(new_n578_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n453_), .A2(new_n510_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(G1336gat));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n508_), .A3(new_n366_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n762_), .A2(new_n366_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n508_), .ZN(G1337gat));
  NAND2_X1  g566(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n413_), .A2(new_n514_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n759_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n762_), .A2(new_n452_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G99gat), .ZN(new_n772_));
  NOR2_X1   g571(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n760_), .A2(new_n535_), .A3(new_n293_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n762_), .A2(new_n293_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(G106gat), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT52), .B(new_n535_), .C1(new_n762_), .C2(new_n293_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g580(.A1(new_n499_), .A2(new_n630_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n673_), .A2(new_n577_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n673_), .A2(new_n577_), .A3(new_n782_), .A4(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n574_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n476_), .A2(new_n481_), .A3(new_n487_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n486_), .A2(new_n479_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n792_), .B(new_n496_), .C1(new_n793_), .C2(new_n487_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n498_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n791_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n567_), .A2(new_n565_), .A3(new_n569_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n570_), .B2(new_n564_), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT55), .B(new_n565_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n505_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n801_), .B2(new_n505_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT58), .B(new_n796_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT115), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n505_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n801_), .A2(KEYINPUT56), .A3(new_n505_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(KEYINPUT58), .A4(new_n796_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n796_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n805_), .A2(new_n812_), .A3(new_n815_), .A4(new_n616_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n795_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n574_), .A2(new_n499_), .A3(KEYINPUT114), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT114), .B1(new_n574_), .B2(new_n499_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n818_), .B1(new_n810_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n817_), .B1(new_n822_), .B2(new_n642_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n820_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n574_), .A2(new_n499_), .A3(KEYINPUT114), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n824_), .B(new_n825_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n818_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n642_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(KEYINPUT57), .A3(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n816_), .A2(new_n823_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n790_), .B1(new_n831_), .B2(new_n630_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n367_), .A2(new_n452_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n832_), .A2(new_n453_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n499_), .B2(KEYINPUT117), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(KEYINPUT117), .B2(new_n837_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n840_));
  OAI211_X1 g639(.A(new_n836_), .B(new_n839_), .C1(new_n834_), .C2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n834_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n837_), .B1(new_n842_), .B2(new_n500_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1340gat));
  XNOR2_X1  g645(.A(KEYINPUT119), .B(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n577_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n834_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n836_), .B(new_n578_), .C1(new_n834_), .C2(new_n840_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n850_), .A2(KEYINPUT120), .ZN(new_n851_));
  INV_X1    g650(.A(new_n847_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n850_), .B2(KEYINPUT120), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n849_), .B1(new_n851_), .B2(new_n853_), .ZN(G1341gat));
  NOR2_X1   g653(.A1(new_n834_), .A2(new_n840_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n727_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G127gat), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n630_), .A2(G127gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n842_), .B2(new_n859_), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n834_), .A2(new_n861_), .A3(new_n642_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n856_), .A2(new_n616_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n861_), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n832_), .A2(new_n453_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n444_), .A2(new_n452_), .A3(new_n366_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n500_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n240_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n577_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n241_), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n867_), .A2(new_n630_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  OAI21_X1  g673(.A(new_n234_), .B1(new_n867_), .B2(new_n829_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n616_), .A2(G162gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT121), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n867_), .B2(new_n877_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT122), .Z(G1347gat));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n414_), .A2(new_n444_), .A3(new_n366_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n500_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n828_), .B2(new_n829_), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n817_), .B(new_n642_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n727_), .B1(new_n885_), .B2(new_n816_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n880_), .B(new_n882_), .C1(new_n886_), .C2(new_n790_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n882_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT123), .B1(new_n832_), .B2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(G169gat), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n887_), .A2(new_n889_), .A3(KEYINPUT124), .A4(G169gat), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n892_), .A2(KEYINPUT62), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n891_), .A3(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n832_), .A2(new_n881_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT22), .B(G169gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n499_), .A2(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT125), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n897_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT126), .B1(new_n894_), .B2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n892_), .A2(KEYINPUT62), .A3(new_n893_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n904_), .A2(new_n896_), .A3(new_n905_), .A4(new_n901_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n906_), .ZN(G1348gat));
  NAND2_X1  g706(.A1(new_n897_), .A2(new_n578_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n897_), .A2(new_n727_), .ZN(new_n910_));
  MUX2_X1   g709(.A(new_n336_), .B(G183gat), .S(new_n910_), .Z(G1350gat));
  NAND4_X1  g710(.A1(new_n897_), .A2(new_n642_), .A3(new_n337_), .A4(new_n302_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n832_), .A2(new_n673_), .A3(new_n881_), .ZN(new_n913_));
  INV_X1    g712(.A(G190gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1351gat));
  NAND4_X1  g714(.A1(new_n453_), .A2(new_n293_), .A3(new_n366_), .A4(new_n413_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n832_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n499_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n578_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n727_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AND2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n922_), .B2(new_n923_), .ZN(G1354gat));
  INV_X1    g725(.A(G218gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n917_), .A2(new_n927_), .A3(new_n642_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n832_), .A2(new_n673_), .A3(new_n916_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n927_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


