//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_;
  INV_X1    g000(.A(G57gat), .ZN(new_n202_));
  INV_X1    g001(.A(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT11), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n210_), .A3(new_n205_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT11), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(KEYINPUT68), .A3(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT6), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT10), .B(G99gat), .Z(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT64), .B(G85gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT9), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G85gat), .ZN(new_n232_));
  INV_X1    g031(.A(G92gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT9), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G85gat), .A2(G92gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n226_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  AND2_X1   g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G85gat), .A2(G92gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(KEYINPUT66), .A3(new_n236_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246_));
  INV_X1    g045(.A(G99gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n225_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n248_), .A2(new_n221_), .A3(new_n222_), .A4(new_n249_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n244_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n245_), .B1(new_n244_), .B2(new_n250_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n238_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n238_), .B(KEYINPUT67), .C1(new_n251_), .C2(new_n252_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n218_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT69), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n218_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n214_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(KEYINPUT12), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT12), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n259_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n259_), .A2(KEYINPUT70), .A3(new_n267_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n257_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n261_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n263_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G120gat), .B(G148gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT72), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT73), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G176gat), .B(G204gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n278_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n263_), .A2(new_n274_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(KEYINPUT13), .ZN(new_n288_));
  XOR2_X1   g087(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n285_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT75), .B(G43gat), .ZN(new_n293_));
  INV_X1    g092(.A(G50gat), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  OR3_X1    g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n297_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT15), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302_));
  INV_X1    g101(.A(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(G8gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT14), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G8gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n300_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n300_), .B(new_n311_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n310_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G113gat), .B(G141gat), .ZN(new_n317_));
  INV_X1    g116(.A(G169gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G197gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n313_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT80), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n292_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n301_), .A2(new_n253_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n255_), .A2(new_n256_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n300_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G232gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT34), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n329_), .B(new_n331_), .C1(KEYINPUT35), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(KEYINPUT35), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G190gat), .B(G218gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G134gat), .ZN(new_n338_));
  INV_X1    g137(.A(G162gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT36), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n334_), .A2(new_n335_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n340_), .B(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n334_), .A2(new_n335_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT37), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G231gat), .A2(G233gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n308_), .B(new_n350_), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(new_n214_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G127gat), .B(G155gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G183gat), .B(G211gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT78), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT79), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n351_), .B(new_n218_), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n357_), .B(KEYINPUT17), .Z(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT37), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n349_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G141gat), .B(G148gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT87), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n372_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT88), .B1(new_n372_), .B2(KEYINPUT1), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI22_X1  g174(.A1(new_n372_), .A2(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n370_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n378_));
  NOR2_X1   g177(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n379_));
  INV_X1    g178(.A(G141gat), .ZN(new_n380_));
  INV_X1    g179(.A(G148gat), .ZN(new_n381_));
  OAI22_X1  g180(.A1(new_n378_), .A2(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n383_));
  OR3_X1    g182(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n386_));
  OAI221_X1 g185(.A(new_n372_), .B1(G155gat), .B2(G162gat), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n377_), .A2(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n388_), .A2(KEYINPUT29), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G78gat), .B(G106gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT28), .Z(new_n394_));
  XNOR2_X1  g193(.A(G211gat), .B(G218gat), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n395_), .A2(KEYINPUT21), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(KEYINPUT21), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G197gat), .B(G204gat), .ZN(new_n398_));
  OR3_X1    g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n395_), .A2(new_n398_), .A3(KEYINPUT21), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n388_), .B2(KEYINPUT29), .ZN(new_n403_));
  INV_X1    g202(.A(G228gat), .ZN(new_n404_));
  INV_X1    g203(.A(G233gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n403_), .A2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n394_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n409_), .A2(new_n394_), .A3(new_n410_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n392_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n411_), .A3(new_n391_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G183gat), .A2(G190gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n421_));
  MUX2_X1   g220(.A(new_n418_), .B(new_n420_), .S(new_n421_), .Z(new_n422_));
  INV_X1    g221(.A(G176gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT24), .B1(new_n318_), .B2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425_));
  MUX2_X1   g224(.A(new_n424_), .B(KEYINPUT24), .S(new_n425_), .Z(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT25), .B(G183gat), .ZN(new_n427_));
  INV_X1    g226(.A(G190gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT81), .B1(new_n428_), .B2(KEYINPUT26), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G190gat), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n427_), .B(new_n429_), .C1(new_n430_), .C2(KEYINPUT81), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n426_), .A3(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n318_), .A2(new_n423_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT22), .B(G169gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n423_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n420_), .A2(KEYINPUT23), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n418_), .A2(new_n421_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(G183gat), .A2(G190gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n435_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n432_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G99gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n443_));
  XNOR2_X1  g242(.A(G15gat), .B(G43gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G71gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n445_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n442_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G127gat), .B(G134gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G113gat), .B(G120gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n456_), .A3(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT31), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT31), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n457_), .A2(new_n462_), .A3(new_n458_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n450_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(new_n464_), .B2(new_n450_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n417_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n459_), .A2(new_n388_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n377_), .A2(new_n455_), .A3(new_n387_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT4), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n459_), .A2(new_n388_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT97), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n478_), .A2(new_n479_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n473_), .B(new_n476_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT98), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n478_), .A2(new_n479_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n480_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT98), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n473_), .A4(new_n476_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n474_), .A2(new_n475_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n472_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n484_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G85gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n484_), .A2(new_n488_), .A3(new_n490_), .A4(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n471_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n427_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n430_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n436_), .A2(new_n437_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(new_n426_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT92), .ZN(new_n507_));
  MUX2_X1   g306(.A(new_n435_), .B(new_n433_), .S(KEYINPUT93), .Z(new_n508_));
  INV_X1    g307(.A(KEYINPUT94), .ZN(new_n509_));
  INV_X1    g308(.A(new_n439_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n508_), .A2(new_n509_), .B1(new_n510_), .B2(new_n422_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n509_), .B2(new_n508_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT20), .B1(new_n441_), .B2(new_n401_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n513_), .A2(new_n401_), .B1(KEYINPUT90), .B2(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n514_), .A2(KEYINPUT90), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G226gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT19), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n441_), .B2(new_n401_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n520_), .B(new_n522_), .C1(new_n513_), .C2(new_n401_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n517_), .A2(new_n519_), .B1(KEYINPUT95), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT18), .B(G64gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(G92gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G8gat), .B(G36gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  OR2_X1    g327(.A1(new_n523_), .A2(KEYINPUT95), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n512_), .A2(new_n402_), .A3(new_n506_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n522_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT102), .B1(new_n532_), .B2(new_n519_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n519_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n535_), .B2(KEYINPUT102), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n530_), .B1(new_n536_), .B2(new_n528_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT27), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n530_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n528_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n538_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT103), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n517_), .A2(new_n519_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n523_), .A2(KEYINPUT95), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n529_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n528_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n530_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(KEYINPUT103), .A3(new_n538_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n539_), .B1(new_n544_), .B2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n501_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n417_), .A2(new_n467_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT33), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n556_), .A2(KEYINPUT100), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n499_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n489_), .A2(new_n473_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n497_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n486_), .A2(new_n476_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n561_), .B2(new_n472_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n550_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(KEYINPUT100), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n499_), .A2(new_n557_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n558_), .A2(new_n563_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT101), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n536_), .B1(new_n567_), .B2(new_n547_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n528_), .A2(KEYINPUT32), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n547_), .A2(KEYINPUT101), .A3(new_n569_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n500_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n555_), .B1(new_n566_), .B2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n328_), .B(new_n369_), .C1(new_n553_), .C2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT104), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT104), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n303_), .A3(new_n500_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT38), .ZN(new_n579_));
  INV_X1    g378(.A(new_n500_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n566_), .A2(new_n572_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n581_), .A2(new_n554_), .B1(new_n501_), .B2(new_n552_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n582_), .A2(new_n327_), .A3(new_n292_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n348_), .B(KEYINPUT105), .Z(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n366_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT106), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT106), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n588_), .A3(new_n585_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n580_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n579_), .B1(new_n303_), .B2(new_n590_), .ZN(G1324gat));
  OAI21_X1  g390(.A(G8gat), .B1(new_n586_), .B2(new_n552_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT39), .ZN(new_n593_));
  AOI21_X1  g392(.A(G8gat), .B1(new_n575_), .B2(new_n576_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n552_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n594_), .A2(KEYINPUT107), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT107), .B1(new_n594_), .B2(new_n595_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n593_), .B(KEYINPUT40), .C1(new_n596_), .C2(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1325gat));
  INV_X1    g401(.A(G15gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n587_), .A2(new_n589_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n467_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(KEYINPUT41), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(KEYINPUT41), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n467_), .A2(new_n603_), .ZN(new_n608_));
  OAI22_X1  g407(.A1(new_n606_), .A2(new_n607_), .B1(new_n574_), .B2(new_n608_), .ZN(G1326gat));
  INV_X1    g408(.A(new_n417_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n611_));
  INV_X1    g410(.A(G22gat), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT42), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(KEYINPUT42), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n417_), .A2(new_n612_), .ZN(new_n616_));
  OAI22_X1  g415(.A1(new_n614_), .A2(new_n615_), .B1(new_n574_), .B2(new_n616_), .ZN(G1327gat));
  INV_X1    g416(.A(new_n348_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n366_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n583_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(G29gat), .B1(new_n622_), .B2(new_n500_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT43), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n349_), .A2(new_n368_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n582_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT43), .B(new_n627_), .C1(new_n553_), .C2(new_n573_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n626_), .A2(new_n628_), .A3(new_n366_), .A4(new_n328_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT44), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(new_n500_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n623_), .B1(new_n631_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g431(.A(G36gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n622_), .A2(new_n633_), .A3(new_n595_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT45), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n630_), .A2(new_n595_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n635_), .B(KEYINPUT46), .C1(new_n636_), .C2(new_n633_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT45), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n634_), .B(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n633_), .B1(new_n630_), .B2(new_n595_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n642_), .ZN(G1329gat));
  AOI21_X1  g442(.A(G43gat), .B1(new_n622_), .B2(new_n467_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n467_), .A2(G43gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n630_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT47), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(G1330gat));
  AOI21_X1  g447(.A(G50gat), .B1(new_n622_), .B2(new_n417_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n610_), .A2(new_n294_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n630_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1331gat));
  NOR2_X1   g452(.A1(new_n582_), .A2(new_n326_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n584_), .A2(new_n366_), .A3(new_n291_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n656_), .A2(new_n202_), .A3(new_n580_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT111), .Z(new_n658_));
  OR3_X1    g457(.A1(new_n582_), .A2(KEYINPUT109), .A3(new_n326_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT109), .B1(new_n582_), .B2(new_n326_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n292_), .A3(new_n369_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n580_), .B1(new_n663_), .B2(KEYINPUT110), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(KEYINPUT110), .B2(new_n663_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n658_), .B1(new_n665_), .B2(new_n202_), .ZN(G1332gat));
  OAI21_X1  g465(.A(G64gat), .B1(new_n656_), .B2(new_n552_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT48), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n595_), .A2(new_n203_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n662_), .B2(new_n669_), .ZN(G1333gat));
  OAI21_X1  g469(.A(G71gat), .B1(new_n656_), .B2(new_n468_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT112), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT49), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n671_), .A2(KEYINPUT112), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n662_), .A2(G71gat), .A3(new_n468_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(G1334gat));
  OAI21_X1  g478(.A(G78gat), .B1(new_n656_), .B2(new_n610_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT50), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n610_), .A2(G78gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n662_), .B2(new_n682_), .ZN(G1335gat));
  AND3_X1   g482(.A1(new_n661_), .A2(new_n292_), .A3(new_n620_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n500_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n626_), .A2(new_n366_), .A3(new_n628_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n500_), .A2(new_n230_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n686_), .A2(new_n327_), .A3(new_n292_), .A4(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n685_), .A2(KEYINPUT113), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT113), .B1(new_n685_), .B2(new_n689_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1336gat));
  AOI21_X1  g491(.A(G92gat), .B1(new_n684_), .B2(new_n595_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n552_), .A2(new_n228_), .A3(new_n227_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n686_), .A2(new_n327_), .A3(new_n292_), .A4(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n693_), .A2(KEYINPUT114), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT114), .B1(new_n693_), .B2(new_n696_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1337gat));
  NAND3_X1  g498(.A1(new_n684_), .A2(new_n224_), .A3(new_n467_), .ZN(new_n700_));
  AND4_X1   g499(.A1(new_n327_), .A2(new_n686_), .A3(new_n292_), .A4(new_n467_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n247_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT51), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT51), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n700_), .B(new_n704_), .C1(new_n247_), .C2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1338gat));
  NAND3_X1  g505(.A1(new_n684_), .A2(new_n225_), .A3(new_n417_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n686_), .A2(new_n327_), .A3(new_n292_), .A4(new_n417_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT52), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G106gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G106gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT53), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT53), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n707_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1339gat));
  NAND3_X1  g515(.A1(new_n369_), .A2(new_n327_), .A3(new_n291_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(KEYINPUT115), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT54), .B1(new_n717_), .B2(KEYINPUT115), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n259_), .A2(KEYINPUT70), .A3(new_n267_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT70), .B1(new_n259_), .B2(new_n267_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n261_), .B(new_n265_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n724_), .B2(new_n257_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n272_), .A2(KEYINPUT55), .A3(new_n261_), .A4(new_n273_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n265_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT69), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n257_), .B(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT116), .B1(new_n728_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n270_), .A2(new_n271_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT116), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n732_), .A2(new_n258_), .A3(new_n733_), .A4(new_n265_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n262_), .A3(new_n734_), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT56), .B(new_n284_), .C1(new_n727_), .C2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(new_n282_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT117), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n326_), .A4(new_n285_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n731_), .A2(new_n262_), .A3(new_n734_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n725_), .A2(new_n726_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n282_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT56), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n738_), .A2(new_n737_), .A3(new_n282_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n746_), .A2(new_n326_), .A3(new_n285_), .A4(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT117), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n314_), .A2(new_n310_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n309_), .A2(new_n312_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT118), .Z(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n752_), .B2(new_n315_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n323_), .B1(new_n753_), .B2(new_n321_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n286_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n742_), .A2(new_n749_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n618_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n746_), .A2(new_n285_), .A3(new_n747_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT120), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(KEYINPUT58), .A4(new_n754_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n746_), .A2(new_n285_), .A3(new_n754_), .A4(new_n747_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT58), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n625_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT120), .B1(new_n764_), .B2(new_n765_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n756_), .A2(KEYINPUT57), .A3(new_n618_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n720_), .B1(new_n770_), .B2(new_n366_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n469_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n595_), .A2(new_n580_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n771_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G113gat), .B1(new_n775_), .B2(new_n326_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n771_), .A2(new_n774_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n469_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NOR4_X1   g579(.A1(new_n771_), .A2(new_n779_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n327_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n776_), .B1(new_n783_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g583(.A(G120gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n291_), .B2(KEYINPUT60), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT121), .Z(new_n787_));
  OAI211_X1 g586(.A(new_n775_), .B(new_n787_), .C1(KEYINPUT60), .C2(new_n785_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n291_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n785_), .ZN(G1341gat));
  AOI21_X1  g589(.A(G127gat), .B1(new_n775_), .B2(new_n619_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n366_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g592(.A(KEYINPUT59), .B1(new_n777_), .B2(new_n469_), .ZN(new_n794_));
  OAI211_X1 g593(.A(G134gat), .B(new_n627_), .C1(new_n794_), .C2(new_n781_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n584_), .ZN(new_n796_));
  NOR4_X1   g595(.A1(new_n771_), .A2(new_n796_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT122), .ZN(new_n798_));
  OR3_X1    g597(.A1(new_n797_), .A2(new_n798_), .A3(G134gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G134gat), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n795_), .A2(new_n799_), .A3(new_n800_), .ZN(G1343gat));
  AOI21_X1  g600(.A(KEYINPUT123), .B1(new_n777_), .B2(new_n470_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n718_), .B(new_n719_), .Z(new_n803_));
  AND3_X1   g602(.A1(new_n756_), .A2(KEYINPUT57), .A3(new_n618_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n758_), .B1(new_n756_), .B2(new_n618_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n763_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n807_), .B2(new_n619_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n808_), .A2(KEYINPUT123), .A3(new_n470_), .A4(new_n773_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n326_), .B1(new_n802_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G141gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n470_), .A3(new_n773_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n809_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(new_n380_), .A3(new_n326_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n817_), .ZN(G1344gat));
  OAI21_X1  g617(.A(new_n292_), .B1(new_n802_), .B2(new_n810_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G148gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n381_), .A3(new_n292_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1345gat));
  XNOR2_X1  g621(.A(KEYINPUT61), .B(G155gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n816_), .B2(new_n619_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n823_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n366_), .B(new_n825_), .C1(new_n815_), .C2(new_n809_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1346gat));
  AOI21_X1  g626(.A(G162gat), .B1(new_n816_), .B2(new_n584_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n339_), .B(new_n625_), .C1(new_n815_), .C2(new_n809_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1347gat));
  NOR2_X1   g629(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n771_), .A2(new_n417_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n552_), .A2(new_n500_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n467_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT124), .Z(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n327_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n318_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n831_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n434_), .ZN(new_n841_));
  OAI221_X1 g640(.A(new_n838_), .B1(KEYINPUT125), .B2(KEYINPUT62), .C1(new_n836_), .C2(new_n327_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(G1348gat));
  NOR2_X1   g642(.A1(new_n836_), .A2(new_n291_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n423_), .ZN(G1349gat));
  AND2_X1   g644(.A1(new_n832_), .A2(new_n835_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n619_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G183gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n503_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1350gat));
  NAND3_X1  g649(.A1(new_n846_), .A2(new_n584_), .A3(new_n430_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G190gat), .B1(new_n836_), .B2(new_n625_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1351gat));
  NAND4_X1  g652(.A1(new_n808_), .A2(new_n326_), .A3(new_n470_), .A4(new_n833_), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n854_), .A2(KEYINPUT126), .A3(new_n320_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n320_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT126), .B1(new_n854_), .B2(new_n320_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(G1352gat));
  AND3_X1   g657(.A1(new_n808_), .A2(new_n470_), .A3(new_n833_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n292_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g660(.A(KEYINPUT63), .B(G211gat), .Z(new_n862_));
  AND3_X1   g661(.A1(new_n859_), .A2(new_n619_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n859_), .A2(new_n619_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1354gat));
  AOI21_X1  g665(.A(G218gat), .B1(new_n859_), .B2(new_n584_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n627_), .A2(G218gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT127), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n859_), .B2(new_n869_), .ZN(G1355gat));
endmodule


