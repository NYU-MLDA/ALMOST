//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_;
  XNOR2_X1  g000(.A(KEYINPUT77), .B(G15gat), .ZN(new_n202_));
  INV_X1    g001(.A(G22gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G1gat), .ZN(new_n205_));
  INV_X1    g004(.A(G8gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G29gat), .B(G36gat), .Z(new_n213_));
  XOR2_X1   g012(.A(G43gat), .B(G50gat), .Z(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT80), .B1(new_n212_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n210_), .A2(new_n218_), .A3(new_n211_), .A4(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n212_), .A2(new_n216_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n222_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G113gat), .B(G141gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G169gat), .B(G197gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n228_), .B(new_n229_), .Z(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT81), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT82), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  OR3_X1    g032(.A1(new_n224_), .A2(new_n227_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n237_));
  XOR2_X1   g036(.A(G85gat), .B(G92gat), .Z(new_n238_));
  NAND2_X1  g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT6), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT6), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(G99gat), .A3(G106gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT64), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  INV_X1    g048(.A(G106gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT65), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(G99gat), .B2(G106gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT7), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n238_), .B1(new_n248_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT8), .B1(new_n238_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  OAI221_X1 g058(.A(new_n238_), .B1(new_n257_), .B2(KEYINPUT8), .C1(new_n248_), .C2(new_n255_), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT10), .B(G99gat), .Z(new_n261_));
  AOI22_X1  g060(.A1(KEYINPUT9), .A2(new_n238_), .B1(new_n261_), .B2(new_n250_), .ZN(new_n262_));
  INV_X1    g061(.A(G85gat), .ZN(new_n263_));
  INV_X1    g062(.A(G92gat), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT9), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n262_), .A2(new_n243_), .A3(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n259_), .A2(new_n260_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G57gat), .B(G64gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G71gat), .B(G78gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(KEYINPUT11), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n272_));
  INV_X1    g071(.A(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n267_), .A2(new_n268_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n259_), .A2(new_n260_), .A3(new_n266_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n259_), .A2(new_n260_), .A3(new_n266_), .A4(new_n276_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT67), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G230gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(KEYINPUT68), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n259_), .A2(new_n260_), .A3(new_n266_), .A4(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n279_), .A2(KEYINPUT12), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT12), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n280_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n281_), .A2(new_n284_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n286_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G120gat), .B(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT5), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G176gat), .B(G204gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT69), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n286_), .A2(new_n296_), .A3(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT13), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n306_), .A2(KEYINPUT13), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n237_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n309_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(KEYINPUT70), .A3(new_n307_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n236_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G228gat), .ZN(new_n314_));
  INV_X1    g113(.A(G233gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G211gat), .B(G218gat), .Z(new_n318_));
  OR2_X1    g117(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n319_));
  INV_X1    g118(.A(G204gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT21), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(G197gat), .B2(G204gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n318_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G197gat), .A2(G204gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n323_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n326_), .A2(new_n327_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n339_));
  AND3_X1   g138(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(KEYINPUT87), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n338_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n335_), .B1(KEYINPUT1), .B2(new_n337_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n337_), .A2(KEYINPUT1), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT29), .B1(new_n348_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n317_), .B1(new_n334_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n334_), .A2(new_n355_), .A3(new_n317_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n358_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n359_), .B1(new_n362_), .B2(new_n356_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(KEYINPUT91), .ZN(new_n366_));
  XOR2_X1   g165(.A(G22gat), .B(G50gat), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT89), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n348_), .A2(new_n354_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NOR4_X1   g171(.A1(new_n348_), .A2(new_n354_), .A3(KEYINPUT89), .A4(KEYINPUT29), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n368_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n342_), .A2(new_n347_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n338_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n354_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n371_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT89), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n370_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n367_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n374_), .A2(new_n375_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n375_), .B1(new_n374_), .B2(new_n383_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n366_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n365_), .A2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n364_), .B(new_n366_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G8gat), .B(G36gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT25), .B(G183gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT26), .B(G190gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT24), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(G169gat), .B2(G176gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n395_), .A2(new_n396_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G183gat), .A2(G190gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT23), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n399_), .A2(new_n397_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n402_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(KEYINPUT92), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n401_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G183gat), .ZN(new_n413_));
  INV_X1    g212(.A(G190gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n405_), .A2(new_n406_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT93), .ZN(new_n417_));
  INV_X1    g216(.A(G169gat), .ZN(new_n418_));
  INV_X1    g217(.A(G176gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT22), .B(G169gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n419_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n405_), .A2(new_n415_), .A3(new_n423_), .A4(new_n406_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n412_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT20), .B1(new_n426_), .B2(new_n334_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT19), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n325_), .A2(new_n328_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n395_), .A2(new_n396_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n398_), .A2(new_n400_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT83), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n401_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n410_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT22), .B1(new_n418_), .B2(KEYINPUT84), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n418_), .A2(KEYINPUT22), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n419_), .B(new_n439_), .C1(new_n440_), .C2(KEYINPUT84), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n441_), .B(new_n416_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n430_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n427_), .A2(new_n429_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n429_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n426_), .B2(new_n334_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n438_), .A2(new_n430_), .A3(new_n442_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n445_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n394_), .B1(new_n444_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n410_), .A2(KEYINPUT92), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n407_), .A2(new_n402_), .A3(new_n408_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n433_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n425_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n334_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n448_), .A2(new_n455_), .A3(KEYINPUT20), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n429_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n453_), .A2(new_n454_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n446_), .B1(new_n458_), .B2(new_n430_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n438_), .A2(new_n442_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n334_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n445_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n394_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n450_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n464_), .A2(KEYINPUT27), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT98), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n429_), .B1(new_n427_), .B2(new_n443_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n447_), .A2(new_n445_), .A3(new_n448_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n472_), .B2(new_n394_), .ZN(new_n473_));
  AOI211_X1 g272(.A(KEYINPUT98), .B(new_n463_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n468_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n389_), .A2(new_n467_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G127gat), .B(G134gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G113gat), .B(G120gat), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G227gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(G15gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G71gat), .B(G99gat), .ZN(new_n485_));
  INV_X1    g284(.A(G43gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n438_), .A2(new_n442_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n488_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n484_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n460_), .A2(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n484_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n489_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n496_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT31), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n492_), .A2(new_n495_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n496_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT31), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n504_), .A2(new_n498_), .A3(new_n505_), .A4(new_n497_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n481_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n477_), .B(new_n478_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n378_), .A2(new_n509_), .A3(new_n379_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n481_), .B1(new_n348_), .B2(new_n354_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G225gat), .A2(G233gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G1gat), .B(G29gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G85gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT0), .B(G57gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT4), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n512_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n511_), .B2(KEYINPUT4), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n513_), .B(new_n518_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT96), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n519_), .B(new_n521_), .C1(KEYINPUT4), .C2(new_n511_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT96), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n513_), .A4(new_n518_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n513_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n517_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n501_), .A2(new_n481_), .A3(new_n506_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n476_), .A2(new_n508_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n463_), .A2(KEYINPUT32), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n444_), .B2(new_n449_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT32), .A4(new_n463_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n530_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT33), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n523_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n510_), .A2(new_n511_), .A3(new_n521_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n517_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT95), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n543_), .A2(new_n546_), .A3(new_n517_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n519_), .B(new_n512_), .C1(KEYINPUT4), .C2(new_n511_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n525_), .A2(KEYINPUT33), .A3(new_n513_), .A4(new_n518_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n542_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n465_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n537_), .A2(new_n530_), .A3(KEYINPUT97), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n540_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n472_), .A2(new_n394_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT98), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n472_), .A2(new_n469_), .A3(new_n394_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n558_), .A2(new_n468_), .B1(new_n466_), .B2(new_n465_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n387_), .A2(new_n531_), .A3(new_n388_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n554_), .A2(new_n389_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n501_), .A2(new_n481_), .A3(new_n506_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(new_n507_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n533_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n313_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT73), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT34), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT71), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n577_), .A2(KEYINPUT71), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n287_), .A2(new_n289_), .A3(new_n225_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n267_), .A2(new_n215_), .B1(new_n576_), .B2(new_n575_), .ZN(new_n583_));
  AOI211_X1 g382(.A(new_n580_), .B(new_n581_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n584_));
  AND4_X1   g383(.A1(KEYINPUT71), .A2(new_n582_), .A3(new_n583_), .A4(new_n577_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n572_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT74), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n583_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n580_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n581_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT71), .A4(new_n577_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT74), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n572_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n593_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n568_), .B(KEYINPUT36), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n587_), .A2(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(KEYINPUT76), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n597_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n594_), .B1(new_n593_), .B2(new_n572_), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT74), .B(new_n571_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n601_), .B(new_n599_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT76), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n597_), .B(KEYINPUT75), .ZN(new_n607_));
  OAI22_X1  g406(.A1(new_n602_), .A2(new_n603_), .B1(new_n593_), .B2(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n600_), .A2(new_n606_), .B1(KEYINPUT37), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n212_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n279_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n610_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n212_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n276_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT79), .B1(new_n612_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617_));
  XOR2_X1   g416(.A(G127gat), .B(G155gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n620_), .B(new_n621_), .Z(new_n622_));
  OR3_X1    g421(.A1(new_n616_), .A2(new_n617_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n625_));
  OAI22_X1  g424(.A1(new_n617_), .A2(new_n625_), .B1(new_n616_), .B2(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n609_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n565_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n205_), .A3(new_n530_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n313_), .A2(new_n627_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n537_), .A2(new_n530_), .A3(KEYINPUT97), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT97), .B1(new_n537_), .B2(new_n530_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n465_), .A2(new_n551_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n389_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n387_), .A2(new_n531_), .A3(new_n388_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n475_), .A2(new_n467_), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n638_), .A2(new_n639_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n508_), .A2(new_n532_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n562_), .A2(new_n507_), .A3(new_n530_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n642_), .A2(new_n643_), .B1(new_n476_), .B2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n598_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n634_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n531_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n631_), .A2(new_n632_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n633_), .A2(new_n649_), .A3(new_n650_), .ZN(G1324gat));
  NAND3_X1  g450(.A1(new_n630_), .A2(new_n206_), .A3(new_n641_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n647_), .A2(new_n641_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  AND4_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .A4(G8gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n206_), .B1(KEYINPUT99), .B2(KEYINPUT39), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n654_), .A2(new_n657_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n652_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1325gat));
  OAI21_X1  g460(.A(G15gat), .B1(new_n648_), .B2(new_n643_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n663_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n630_), .A2(new_n483_), .A3(new_n563_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .ZN(G1326gat));
  AOI21_X1  g466(.A(new_n203_), .B1(new_n647_), .B2(new_n639_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT42), .Z(new_n669_));
  NAND3_X1  g468(.A1(new_n630_), .A2(new_n203_), .A3(new_n639_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1327gat));
  INV_X1    g470(.A(new_n598_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n627_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n565_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n530_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n609_), .A2(new_n564_), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n609_), .B2(new_n564_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n628_), .B(new_n313_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n313_), .A2(new_n628_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n608_), .A2(KEYINPUT37), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT76), .B1(new_n598_), .B2(new_n599_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n604_), .A2(new_n605_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n645_), .B2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n609_), .A2(new_n564_), .A3(new_n676_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n683_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n682_), .B1(new_n690_), .B2(KEYINPUT44), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n679_), .A2(KEYINPUT101), .A3(new_n680_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n681_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n530_), .A2(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n675_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n693_), .B2(new_n641_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n559_), .A2(G36gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n565_), .A2(new_n673_), .A3(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT102), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT102), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n701_), .A2(KEYINPUT45), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n696_), .B1(new_n698_), .B2(new_n707_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n701_), .A2(KEYINPUT45), .A3(new_n702_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT45), .B1(new_n701_), .B2(new_n702_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n559_), .B(new_n681_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n711_), .B(KEYINPUT46), .C1(new_n712_), .C2(new_n697_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n708_), .A2(new_n713_), .ZN(G1329gat));
  AOI21_X1  g513(.A(G43gat), .B1(new_n674_), .B2(new_n563_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n643_), .A2(new_n486_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n693_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(G1330gat));
  INV_X1    g518(.A(G50gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n674_), .A2(new_n720_), .A3(new_n639_), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT103), .B(new_n720_), .C1(new_n693_), .C2(new_n639_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n691_), .A2(new_n692_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n681_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n639_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n723_), .B1(new_n726_), .B2(G50gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n721_), .B1(new_n722_), .B2(new_n727_), .ZN(G1331gat));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729_));
  INV_X1    g528(.A(new_n236_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT105), .B1(new_n645_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n564_), .A2(new_n732_), .A3(new_n236_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n310_), .A2(new_n312_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n609_), .A2(new_n735_), .A3(new_n628_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT104), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(KEYINPUT104), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n729_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n739_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n741_), .A2(KEYINPUT106), .A3(new_n734_), .A4(new_n737_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n531_), .A2(G57gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n627_), .A2(new_n236_), .ZN(new_n745_));
  NOR4_X1   g544(.A1(new_n645_), .A2(new_n735_), .A3(new_n598_), .A4(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G57gat), .B1(new_n747_), .B2(new_n531_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT107), .ZN(G1332gat));
  INV_X1    g549(.A(G64gat), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n740_), .A2(new_n742_), .A3(new_n751_), .A4(new_n641_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n746_), .B2(new_n641_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT109), .ZN(G1333gat));
  INV_X1    g556(.A(G71gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n746_), .B2(new_n563_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT49), .Z(new_n760_));
  NAND4_X1  g559(.A1(new_n740_), .A2(new_n742_), .A3(new_n758_), .A4(new_n563_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1334gat));
  OAI21_X1  g563(.A(G78gat), .B1(new_n747_), .B2(new_n389_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n389_), .A2(G78gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n740_), .A2(new_n742_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1335gat));
  NOR3_X1   g569(.A1(new_n735_), .A2(new_n627_), .A3(new_n672_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n734_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n263_), .A3(new_n530_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n688_), .A2(new_n689_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n735_), .A2(new_n627_), .A3(new_n730_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(new_n530_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n777_), .B2(new_n263_), .ZN(G1336gat));
  AOI21_X1  g577(.A(new_n264_), .B1(new_n776_), .B2(new_n641_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n559_), .A2(G92gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT112), .ZN(G1337gat));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n563_), .A2(new_n261_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n636_), .A2(new_n637_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n639_), .B1(new_n785_), .B2(new_n553_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n641_), .A2(new_n640_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n643_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT105), .B(new_n730_), .C1(new_n788_), .C2(new_n533_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n732_), .B1(new_n564_), .B2(new_n236_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n771_), .B(new_n784_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n734_), .A2(KEYINPUT113), .A3(new_n771_), .A4(new_n784_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n563_), .B(new_n775_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n793_), .A2(new_n794_), .B1(G99gat), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n783_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT51), .B1(new_n796_), .B2(KEYINPUT114), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n793_), .A2(new_n794_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n795_), .A2(G99gat), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(KEYINPUT114), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n801_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n796_), .A2(KEYINPUT114), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n806_), .A2(new_n783_), .A3(new_n807_), .A4(KEYINPUT51), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n803_), .A2(new_n808_), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n772_), .A2(new_n250_), .A3(new_n639_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n774_), .A2(new_n639_), .A3(new_n775_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(G106gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(G106gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI211_X1 g615(.A(new_n627_), .B(new_n236_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n609_), .A2(KEYINPUT54), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n308_), .A2(new_n309_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n745_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n687_), .B2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  INV_X1    g623(.A(new_n230_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n221_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n230_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n304_), .A2(new_n305_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n234_), .A2(new_n235_), .A3(new_n305_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n296_), .A2(KEYINPUT55), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n292_), .A2(new_n294_), .A3(new_n835_), .A4(new_n295_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n292_), .A2(new_n294_), .A3(new_n282_), .A4(new_n277_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n834_), .A2(new_n836_), .B1(new_n285_), .B2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n302_), .B1(new_n838_), .B2(KEYINPUT116), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n285_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT117), .B1(new_n839_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n833_), .B1(new_n845_), .B2(KEYINPUT56), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n840_), .A2(KEYINPUT116), .A3(new_n841_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n303_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n838_), .A2(KEYINPUT116), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n832_), .B1(new_n846_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n824_), .B1(new_n854_), .B2(new_n598_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n847_), .B(KEYINPUT56), .C1(new_n849_), .C2(new_n850_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n234_), .A2(new_n235_), .A3(new_n305_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n839_), .A2(new_n844_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT56), .B1(new_n859_), .B2(new_n847_), .ZN(new_n860_));
  OAI22_X1  g659(.A1(new_n858_), .A2(new_n860_), .B1(new_n831_), .B2(new_n830_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(KEYINPUT57), .A3(new_n672_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(KEYINPUT56), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n839_), .A2(new_n844_), .A3(new_n852_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n828_), .A2(new_n829_), .A3(new_n305_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n863_), .A2(KEYINPUT58), .A3(new_n864_), .A4(new_n865_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n609_), .A3(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n855_), .A2(new_n862_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n823_), .B1(new_n628_), .B2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n563_), .A2(new_n530_), .A3(new_n476_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G113gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n730_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n871_), .A2(new_n628_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n823_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n873_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(KEYINPUT59), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n236_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n876_), .B1(new_n884_), .B2(new_n875_), .ZN(G1340gat));
  INV_X1    g684(.A(G120gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n735_), .B2(KEYINPUT60), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n874_), .B(new_n887_), .C1(KEYINPUT60), .C2(new_n886_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n735_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n886_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n874_), .A2(new_n891_), .A3(new_n627_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n628_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1342gat));
  INV_X1    g693(.A(G134gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n687_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT59), .B1(new_n879_), .B2(new_n880_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n872_), .A2(new_n882_), .A3(new_n873_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n874_), .A2(new_n598_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n895_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n899_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n896_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G134gat), .B1(new_n874_), .B2(new_n598_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT118), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n907_), .ZN(G1343gat));
  NOR4_X1   g707(.A1(new_n563_), .A2(new_n531_), .A3(new_n389_), .A4(new_n641_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n872_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n730_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g712(.A(new_n735_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g715(.A1(new_n879_), .A2(new_n909_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT119), .B1(new_n917_), .B2(new_n628_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n911_), .A2(new_n919_), .A3(new_n627_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n918_), .A2(new_n920_), .A3(new_n922_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1346gat));
  OR3_X1    g725(.A1(new_n917_), .A2(G162gat), .A3(new_n672_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G162gat), .B1(new_n917_), .B2(new_n687_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1347gat));
  NAND2_X1  g728(.A1(new_n644_), .A2(new_n641_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n872_), .A2(new_n639_), .A3(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n931_), .A2(new_n421_), .A3(new_n730_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n639_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n930_), .A2(new_n236_), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n935_), .B(KEYINPUT120), .Z(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n933_), .B1(new_n937_), .B2(G169gat), .ZN(new_n938_));
  AOI211_X1 g737(.A(KEYINPUT62), .B(new_n418_), .C1(new_n934_), .C2(new_n936_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n932_), .B1(new_n938_), .B2(new_n939_), .ZN(G1348gat));
  NAND2_X1  g739(.A1(new_n931_), .A2(new_n914_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(KEYINPUT121), .A2(G176gat), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(KEYINPUT121), .B(G176gat), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n941_), .B2(new_n944_), .ZN(G1349gat));
  INV_X1    g744(.A(new_n930_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n879_), .A2(new_n627_), .A3(new_n389_), .A4(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n413_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n949_));
  INV_X1    g748(.A(new_n395_), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n934_), .A2(new_n627_), .A3(new_n950_), .A4(new_n946_), .ZN(new_n951_));
  AND3_X1   g750(.A1(new_n948_), .A2(new_n949_), .A3(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n949_), .B1(new_n948_), .B2(new_n951_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n931_), .A2(new_n598_), .A3(new_n396_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n931_), .A2(new_n609_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n414_), .ZN(G1351gat));
  XOR2_X1   g756(.A(KEYINPUT123), .B(G197gat), .Z(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT123), .A2(G197gat), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n563_), .A2(new_n640_), .A3(new_n559_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n879_), .A2(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n236_), .ZN(new_n962_));
  MUX2_X1   g761(.A(new_n958_), .B(new_n959_), .S(new_n962_), .Z(G1352gat));
  NOR2_X1   g762(.A1(new_n961_), .A2(new_n735_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(new_n320_), .ZN(G1353gat));
  INV_X1    g764(.A(new_n961_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n627_), .A2(new_n967_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(KEYINPUT124), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n969_), .B1(KEYINPUT125), .B2(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n966_), .A2(new_n971_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n970_), .A2(KEYINPUT125), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n972_), .B(new_n973_), .ZN(G1354gat));
  XOR2_X1   g773(.A(KEYINPUT126), .B(G218gat), .Z(new_n975_));
  NOR3_X1   g774(.A1(new_n961_), .A2(new_n687_), .A3(new_n975_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n966_), .A2(new_n598_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n975_), .ZN(G1355gat));
endmodule


