//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT3), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  AND2_X1   g003(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n203_), .B(new_n207_), .C1(new_n204_), .C2(new_n206_), .ZN(new_n208_));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n202_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT87), .ZN(new_n218_));
  INV_X1    g017(.A(new_n210_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n209_), .B2(new_n216_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n204_), .B(new_n215_), .C1(new_n218_), .C2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G197gat), .B(G204gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n225_), .A2(KEYINPUT21), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n226_), .B(KEYINPUT93), .Z(new_n227_));
  INV_X1    g026(.A(G204gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n229_));
  OAI211_X1 g028(.A(KEYINPUT21), .B(new_n229_), .C1(new_n225_), .C2(KEYINPUT91), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G211gat), .B(G218gat), .Z(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n227_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n225_), .A2(KEYINPUT21), .A3(new_n233_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n223_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G78gat), .B(G106gat), .Z(new_n242_));
  OAI21_X1  g041(.A(new_n223_), .B1(KEYINPUT90), .B2(new_n240_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(KEYINPUT90), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n235_), .A2(KEYINPUT94), .A3(new_n236_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT94), .B1(new_n235_), .B2(new_n236_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n241_), .B(new_n242_), .C1(new_n243_), .C2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT95), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G22gat), .B(G50gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT28), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n250_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n241_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n242_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n248_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n249_), .A2(new_n248_), .A3(new_n257_), .A4(new_n253_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G8gat), .B(G36gat), .ZN(new_n262_));
  INV_X1    g061(.A(G92gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT18), .B(G64gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT84), .B(G176gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT22), .B(G169gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT85), .ZN(new_n272_));
  INV_X1    g071(.A(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT23), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G183gat), .A3(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(G183gat), .B2(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n272_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n277_), .B(KEYINPUT83), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n275_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n267_), .A2(KEYINPUT24), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  MUX2_X1   g083(.A(new_n283_), .B(KEYINPUT24), .S(new_n284_), .Z(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G190gat), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n273_), .A2(KEYINPUT25), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n273_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT82), .B1(new_n273_), .B2(KEYINPUT25), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n286_), .B(new_n287_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n282_), .A2(new_n285_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n282_), .B1(G183gat), .B2(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n269_), .A2(new_n270_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n267_), .B(KEYINPUT98), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT25), .B(G183gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n286_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n285_), .A2(new_n278_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT20), .B1(new_n237_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n293_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n306_), .B(KEYINPUT97), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n246_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n235_), .A2(KEYINPUT94), .A3(new_n236_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n292_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT20), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n237_), .B2(new_n301_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n310_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n266_), .B1(new_n308_), .B2(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n245_), .A2(new_n246_), .A3(new_n292_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n316_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n309_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n293_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n266_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(KEYINPUT99), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT99), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n321_), .A2(new_n326_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G85gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT0), .B(G57gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  XNOR2_X1  g131(.A(G127gat), .B(G134gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G113gat), .B(G120gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n222_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n214_), .A2(new_n221_), .A3(new_n335_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(KEYINPUT4), .A3(new_n338_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n222_), .A2(new_n344_), .A3(new_n336_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n340_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n332_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT100), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT100), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n349_), .B(new_n332_), .C1(new_n342_), .C2(new_n346_), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT101), .B(KEYINPUT33), .Z(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  OAI211_X1 g151(.A(KEYINPUT33), .B(new_n332_), .C1(new_n342_), .C2(new_n346_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT102), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n343_), .A2(new_n345_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n341_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n332_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n343_), .A2(KEYINPUT102), .A3(new_n340_), .A4(new_n345_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n328_), .A2(new_n352_), .A3(new_n353_), .A4(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n339_), .A2(new_n341_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n341_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n332_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n347_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n323_), .A2(KEYINPUT32), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n321_), .A2(new_n322_), .A3(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n319_), .A2(new_n320_), .A3(new_n309_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n302_), .A2(KEYINPUT103), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n302_), .A2(KEYINPUT103), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n293_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n371_), .B2(new_n306_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n365_), .B(new_n367_), .C1(new_n372_), .C2(new_n366_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n261_), .B1(new_n360_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G71gat), .B(G99gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G227gat), .ZN(new_n377_));
  INV_X1    g176(.A(G233gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n313_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n280_), .B2(new_n291_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n292_), .A2(KEYINPUT30), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n386_), .A2(new_n379_), .A3(new_n383_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G15gat), .B(G43gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n382_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n379_), .B1(new_n386_), .B2(new_n383_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n335_), .B(KEYINPUT31), .Z(new_n394_));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n390_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n389_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(new_n392_), .A3(new_n388_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n376_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n396_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n400_), .A3(new_n398_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n375_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n260_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n249_), .A2(new_n253_), .B1(new_n257_), .B2(new_n248_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n405_), .B(new_n402_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n260_), .A3(new_n259_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT104), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n365_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n364_), .A2(new_n347_), .A3(KEYINPUT104), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT27), .B(new_n324_), .C1(new_n372_), .C2(new_n323_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT27), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n325_), .A2(new_n418_), .A3(new_n327_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n374_), .A2(new_n407_), .B1(new_n412_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G230gat), .A2(G233gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n422_), .B(KEYINPUT64), .Z(new_n423_));
  XNOR2_X1  g222(.A(G57gat), .B(G64gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT11), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G71gat), .B(G78gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n425_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n424_), .A2(KEYINPUT11), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n427_), .B1(new_n430_), .B2(new_n426_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G99gat), .A2(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT6), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(G99gat), .A3(G106gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n438_));
  INV_X1    g237(.A(G99gat), .ZN(new_n439_));
  INV_X1    g238(.A(G106gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT7), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT67), .B1(G99gat), .B2(G106gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n445_), .A2(KEYINPUT68), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n441_), .A2(new_n448_), .A3(new_n442_), .A4(new_n443_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n437_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G85gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(new_n263_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT8), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n447_), .A2(new_n449_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT70), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT69), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT70), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n436_), .B(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n454_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n457_), .B1(new_n465_), .B2(KEYINPUT8), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT10), .B(G99gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n437_), .B1(new_n440_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT9), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT65), .B(G92gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(new_n451_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT66), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n453_), .B1(new_n452_), .B2(KEYINPUT9), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n470_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n431_), .B1(new_n466_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n454_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n436_), .A2(new_n463_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n433_), .A2(new_n435_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n447_), .A2(new_n449_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n483_), .A2(new_n455_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n431_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n473_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n475_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n469_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n477_), .A2(KEYINPUT12), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n489_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT12), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n431_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n423_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n423_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n477_), .B2(new_n490_), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n498_));
  XNOR2_X1  g297(.A(G120gat), .B(G148gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G176gat), .B(G204gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n495_), .A2(new_n497_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n507_), .A2(KEYINPUT13), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(KEYINPUT13), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT81), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512_));
  INV_X1    g311(.A(G1gat), .ZN(new_n513_));
  INV_X1    g312(.A(G8gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G8gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G29gat), .B(G36gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT78), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n521_), .B(KEYINPUT15), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n518_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT79), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n518_), .A2(new_n522_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n524_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(G229gat), .A3(G233gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G169gat), .B(G197gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n534_), .A2(KEYINPUT80), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n534_), .B2(KEYINPUT80), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n511_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(KEYINPUT81), .A3(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n421_), .A2(new_n510_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT34), .Z(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n525_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT73), .ZN(new_n556_));
  OAI22_X1  g355(.A1(new_n555_), .A2(new_n556_), .B1(new_n492_), .B2(new_n522_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n492_), .A2(new_n525_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(KEYINPUT73), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n553_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n550_), .B(new_n551_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n558_), .B(new_n561_), .C1(new_n492_), .C2(new_n522_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT36), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT74), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n566_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(KEYINPUT36), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n560_), .A2(new_n572_), .A3(new_n562_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n548_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT75), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n568_), .B1(new_n563_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n560_), .A2(KEYINPUT75), .A3(new_n562_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n575_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n580_));
  AOI21_X1  g379(.A(new_n574_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n518_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(new_n431_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G211gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT16), .B(G183gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT77), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n584_), .A2(new_n591_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(KEYINPUT17), .B2(new_n588_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n581_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n547_), .A2(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n599_), .A2(G1gat), .A3(new_n416_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT38), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n421_), .A2(new_n579_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n540_), .A2(new_n541_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n510_), .A2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n602_), .A2(new_n596_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n416_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n600_), .A2(KEYINPUT38), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n601_), .A2(new_n608_), .A3(new_n609_), .ZN(G1324gat));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n419_), .A2(new_n417_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n606_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n611_), .B1(new_n614_), .B2(G8gat), .ZN(new_n615_));
  AOI211_X1 g414(.A(KEYINPUT39), .B(new_n514_), .C1(new_n606_), .C2(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n514_), .ZN(new_n617_));
  OAI22_X1  g416(.A1(new_n615_), .A2(new_n616_), .B1(new_n599_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n607_), .B2(new_n407_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT105), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT41), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n599_), .A2(G15gat), .A3(new_n407_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n621_), .A2(KEYINPUT105), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(KEYINPUT105), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT41), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n625_), .A3(new_n628_), .ZN(G1326gat));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n606_), .B2(new_n261_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT42), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n261_), .A2(new_n630_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n599_), .B2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(new_n581_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT43), .B1(new_n421_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n261_), .B(new_n406_), .C1(new_n360_), .C2(new_n373_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n637_), .B(new_n581_), .C1(new_n638_), .C2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n605_), .A2(new_n597_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT106), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n416_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n642_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G29gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n579_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n596_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n547_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n416_), .A2(G29gat), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT107), .Z(new_n658_));
  OAI21_X1  g457(.A(new_n652_), .B1(new_n656_), .B2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(G36gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n655_), .A2(new_n660_), .A3(new_n613_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n662_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n655_), .A2(new_n660_), .A3(new_n613_), .A4(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n612_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n660_), .B1(new_n667_), .B2(new_n650_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n666_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1329gat));
  NAND4_X1  g471(.A1(new_n648_), .A2(G43gat), .A3(new_n406_), .A4(new_n650_), .ZN(new_n673_));
  INV_X1    g472(.A(G43gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n656_), .B2(new_n407_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g476(.A(G50gat), .B1(new_n655_), .B2(new_n261_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n648_), .A2(new_n261_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n650_), .A2(G50gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(G1331gat));
  INV_X1    g480(.A(G57gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n510_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n603_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n421_), .A2(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(new_n598_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT109), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n649_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n687_), .A2(KEYINPUT109), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n682_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n692_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n542_), .A2(new_n544_), .A3(new_n596_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n602_), .A2(new_n510_), .A3(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT111), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT112), .B(G57gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n416_), .A2(new_n698_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n693_), .A2(new_n694_), .B1(new_n697_), .B2(new_n699_), .ZN(G1332gat));
  INV_X1    g499(.A(G64gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n687_), .A2(new_n701_), .A3(new_n613_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n697_), .A2(new_n613_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(G64gat), .ZN(new_n705_));
  AOI211_X1 g504(.A(KEYINPUT48), .B(new_n701_), .C1(new_n697_), .C2(new_n613_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1333gat));
  INV_X1    g506(.A(G71gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n687_), .A2(new_n708_), .A3(new_n406_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n697_), .A2(new_n406_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(G71gat), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT49), .B(new_n708_), .C1(new_n697_), .C2(new_n406_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(G1334gat));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n687_), .A2(new_n715_), .A3(new_n261_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT50), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n697_), .A2(new_n261_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G78gat), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT50), .B(new_n715_), .C1(new_n697_), .C2(new_n261_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1335gat));
  AND2_X1   g520(.A1(new_n686_), .A2(new_n654_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n649_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT113), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n596_), .B(new_n685_), .C1(new_n636_), .C2(new_n641_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n416_), .A2(new_n451_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n722_), .B2(new_n613_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n612_), .A2(new_n472_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n725_), .B2(new_n729_), .ZN(G1337gat));
  NAND4_X1  g529(.A1(new_n642_), .A2(new_n597_), .A3(new_n406_), .A4(new_n684_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n731_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT114), .B1(new_n731_), .B2(G99gat), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n722_), .A2(new_n468_), .A3(new_n406_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n734_), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n731_), .A2(G99gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n731_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n735_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n742_));
  OR2_X1    g541(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n736_), .A2(new_n744_), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n722_), .A2(new_n440_), .A3(new_n261_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n642_), .A2(new_n597_), .A3(new_n261_), .A4(new_n684_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(G106gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G106gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g551(.A(new_n695_), .B1(new_n509_), .B2(new_n508_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT116), .B1(new_n753_), .B2(new_n581_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n683_), .A2(new_n635_), .A3(new_n755_), .A4(new_n695_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(KEYINPUT54), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT116), .B(new_n758_), .C1(new_n753_), .C2(new_n581_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT56), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n491_), .A2(new_n494_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT55), .B1(new_n762_), .B2(new_n496_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n764_), .B(new_n423_), .C1(new_n491_), .C2(new_n494_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n491_), .A2(new_n423_), .A3(new_n494_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n763_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT117), .B(new_n761_), .C1(new_n768_), .C2(new_n502_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n496_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n764_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n495_), .A2(KEYINPUT55), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n766_), .A3(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n503_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n769_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n503_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT117), .B1(new_n776_), .B2(new_n761_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n505_), .B(new_n603_), .C1(new_n775_), .C2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n527_), .A2(new_n529_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n524_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n537_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n530_), .A2(new_n533_), .A3(new_n538_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n507_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n778_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n653_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(KEYINPUT57), .A3(new_n653_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n783_), .A2(new_n505_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n761_), .B1(new_n768_), .B2(new_n502_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n774_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n581_), .B1(new_n792_), .B2(KEYINPUT58), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(KEYINPUT58), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n581_), .B(KEYINPUT118), .C1(new_n792_), .C2(KEYINPUT58), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n788_), .A2(new_n789_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n760_), .B1(new_n799_), .B2(new_n597_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n613_), .A2(new_n416_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n411_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n800_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G113gat), .B1(new_n804_), .B2(new_n603_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n760_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n785_), .B2(new_n653_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n787_), .B(new_n579_), .C1(new_n778_), .C2(new_n784_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n810_), .B2(new_n596_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n803_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT120), .B1(new_n813_), .B2(KEYINPUT59), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n812_), .B2(KEYINPUT120), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n800_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n546_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n805_), .B1(new_n820_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g620(.A(new_n818_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT59), .B1(new_n811_), .B2(new_n822_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n800_), .A2(new_n803_), .A3(new_n814_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n510_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT121), .B(G120gat), .Z(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT122), .B(new_n510_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n828_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n804_), .B(new_n832_), .C1(KEYINPUT60), .C2(new_n831_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(G1341gat));
  AOI21_X1  g633(.A(G127gat), .B1(new_n804_), .B2(new_n596_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n597_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g636(.A(G134gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n804_), .A2(new_n838_), .A3(new_n579_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n635_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT123), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n843_), .B(new_n839_), .C1(new_n840_), .C2(new_n838_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1343gat));
  NOR2_X1   g644(.A1(new_n800_), .A2(new_n410_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n801_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n604_), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n683_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(G148gat), .Z(G1345gat));
  NAND3_X1  g650(.A1(new_n846_), .A2(new_n596_), .A3(new_n801_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT124), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n846_), .A2(new_n854_), .A3(new_n596_), .A4(new_n801_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n853_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1346gat));
  INV_X1    g658(.A(G162gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n847_), .A2(new_n860_), .A3(new_n635_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n847_), .B2(new_n653_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT125), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n864_), .B(new_n860_), .C1(new_n847_), .C2(new_n653_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n861_), .B1(new_n863_), .B2(new_n865_), .ZN(G1347gat));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n612_), .A2(new_n649_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n811_), .A2(new_n802_), .A3(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n604_), .ZN(new_n870_));
  INV_X1    g669(.A(G169gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n270_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT62), .B(G169gat), .C1(new_n869_), .C2(new_n604_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(G1348gat));
  INV_X1    g674(.A(new_n869_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n510_), .ZN(new_n877_));
  INV_X1    g676(.A(G176gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n269_), .B2(new_n877_), .ZN(G1349gat));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n596_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n298_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n273_), .B2(new_n881_), .ZN(G1350gat));
  NAND3_X1  g682(.A1(new_n876_), .A2(new_n579_), .A3(new_n286_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G190gat), .B1(new_n869_), .B2(new_n635_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1351gat));
  NAND2_X1  g685(.A1(new_n846_), .A2(new_n868_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n603_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g689(.A1(new_n887_), .A2(new_n683_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n228_), .ZN(G1353gat));
  NOR2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  AND2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n887_), .A2(new_n597_), .A3(new_n893_), .A4(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n887_), .B2(new_n597_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(KEYINPUT126), .B(new_n893_), .C1(new_n887_), .C2(new_n597_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n895_), .B1(new_n898_), .B2(new_n899_), .ZN(G1354gat));
  AND3_X1   g699(.A1(new_n888_), .A2(G218gat), .A3(new_n581_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G218gat), .B1(new_n888_), .B2(new_n579_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1355gat));
endmodule


