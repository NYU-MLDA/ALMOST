//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT67), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n202_), .A2(new_n203_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G85gat), .B(G92gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT64), .Z(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT6), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT65), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT7), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n214_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n216_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n221_), .ZN(new_n223_));
  OAI22_X1  g022(.A1(new_n220_), .A2(new_n221_), .B1(new_n214_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT9), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n213_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT10), .B(G99gat), .Z(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(G85gat), .A3(G92gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n226_), .A2(new_n229_), .A3(new_n216_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT66), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n224_), .A2(new_n234_), .A3(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n212_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT12), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n212_), .A2(new_n237_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G230gat), .A2(G233gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n210_), .A2(KEYINPUT12), .A3(new_n232_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n212_), .B2(new_n237_), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n245_), .B(new_n240_), .Z(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n246_), .B2(new_n242_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G120gat), .B(G148gat), .ZN(new_n248_));
  INV_X1    g047(.A(G204gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT5), .ZN(new_n251_));
  INV_X1    g050(.A(G176gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n247_), .B(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n255_), .A2(KEYINPUT13), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(KEYINPUT13), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT70), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT74), .B(G1gat), .Z(new_n261_));
  INV_X1    g060(.A(G8gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT14), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G15gat), .B(G22gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G1gat), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n266_), .A2(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n262_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G29gat), .B(G36gat), .ZN(new_n270_));
  INV_X1    g069(.A(G43gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G50gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT77), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n269_), .B(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G229gat), .A3(G233gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT78), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n274_), .B(KEYINPUT15), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n279_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G229gat), .A2(G233gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT79), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G113gat), .B(G141gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(G197gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT80), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n278_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(KEYINPUT24), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT25), .B(G183gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n296_), .A2(KEYINPUT24), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308_));
  NAND3_X1  g107(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(KEYINPUT23), .ZN(new_n311_));
  AOI22_X1  g110(.A1(KEYINPUT81), .A2(new_n304_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n302_), .B(new_n312_), .C1(KEYINPUT81), .C2(new_n304_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(KEYINPUT23), .A3(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n308_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n314_), .B(new_n315_), .C1(G183gat), .C2(G190gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n303_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT22), .B(G169gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(new_n252_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n313_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT83), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G71gat), .B(G99gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G15gat), .B(G43gat), .Z(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT30), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n326_), .B(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n329_), .A2(KEYINPUT84), .ZN(new_n330_));
  XOR2_X1   g129(.A(G127gat), .B(G134gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G113gat), .ZN(new_n332_));
  INV_X1    g131(.A(G120gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT31), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n330_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G22gat), .B(G50gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT86), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n343_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n345_), .A3(KEYINPUT1), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G141gat), .ZN(new_n351_));
  INV_X1    g150(.A(G148gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n347_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT87), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n351_), .B(new_n352_), .C1(KEYINPUT87), .C2(KEYINPUT3), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n355_), .B(new_n356_), .C1(G141gat), .C2(G148gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT88), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n363_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT89), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n340_), .A2(new_n343_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n369_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n354_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT90), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT90), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n376_), .B(new_n354_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT91), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n374_), .A2(KEYINPUT91), .A3(new_n375_), .A4(new_n377_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n338_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(new_n383_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n381_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n337_), .A3(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G78gat), .B(G106gat), .Z(new_n391_));
  OR2_X1    g190(.A1(new_n391_), .A2(KEYINPUT98), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n386_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n368_), .A2(new_n370_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT89), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n376_), .B1(new_n398_), .B2(new_n354_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n377_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT29), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402_));
  OR2_X1    g201(.A1(KEYINPUT93), .A2(G197gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(KEYINPUT93), .A2(G197gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n249_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT94), .ZN(new_n406_));
  INV_X1    g205(.A(G197gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G204gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n403_), .A2(new_n409_), .A3(new_n249_), .A4(new_n404_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT21), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT95), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n249_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n407_), .A2(G204gat), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n414_), .A2(KEYINPUT21), .A3(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(G211gat), .A2(G218gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G211gat), .A2(G218gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n411_), .A2(new_n420_), .A3(KEYINPUT21), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n413_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n418_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT96), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT21), .B1(new_n414_), .B2(new_n415_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT97), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n426_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n423_), .B(KEYINPUT96), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n422_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n401_), .A2(new_n402_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT99), .ZN(new_n435_));
  INV_X1    g234(.A(new_n373_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n433_), .B1(new_n436_), .B2(new_n375_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(G228gat), .A3(G233gat), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n434_), .A2(new_n435_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n435_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n393_), .A2(new_n394_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n391_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n384_), .A2(new_n385_), .A3(new_n338_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n337_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n386_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n443_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n442_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n334_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT102), .B1(new_n452_), .B2(KEYINPUT4), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n451_), .A2(new_n373_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(KEYINPUT4), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n334_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT102), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n453_), .A2(new_n456_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G225gat), .A2(G233gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n463_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT0), .B(G57gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(G85gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(G1gat), .B(G29gat), .Z(new_n471_));
  XOR2_X1   g270(.A(new_n470_), .B(new_n471_), .Z(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n465_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT33), .B1(new_n475_), .B2(new_n472_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n453_), .A2(new_n456_), .A3(new_n462_), .A4(new_n460_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT103), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n452_), .A2(new_n479_), .A3(new_n455_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT103), .B1(new_n457_), .B2(new_n454_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n463_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n472_), .A3(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT18), .B(G64gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G92gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G8gat), .B(G36gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  AND3_X1   g286(.A1(new_n304_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n310_), .A2(new_n311_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n489_), .B1(G183gat), .B2(G190gat), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n302_), .A2(new_n488_), .B1(new_n490_), .B2(new_n319_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT20), .B1(new_n433_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G226gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT100), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT19), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n433_), .A2(new_n321_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n500_));
  INV_X1    g299(.A(new_n433_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n321_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT101), .B1(new_n433_), .B2(new_n492_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT101), .ZN(new_n506_));
  AOI211_X1 g305(.A(new_n506_), .B(new_n491_), .C1(new_n422_), .C2(new_n432_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n503_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n487_), .B(new_n499_), .C1(new_n509_), .C2(new_n497_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n487_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n504_), .A2(new_n507_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n497_), .B1(new_n512_), .B2(new_n503_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n494_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n483_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT104), .B1(new_n477_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT104), .ZN(new_n519_));
  AOI211_X1 g318(.A(new_n519_), .B(new_n516_), .C1(new_n474_), .C2(new_n476_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n467_), .A2(new_n473_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n475_), .A2(new_n472_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n487_), .A2(KEYINPUT32), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n499_), .B(new_n526_), .C1(new_n509_), .C2(new_n497_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n493_), .A2(KEYINPUT105), .B1(new_n433_), .B2(new_n321_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT105), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n529_), .B(KEYINPUT20), .C1(new_n433_), .C2(new_n492_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n497_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  AND4_X1   g330(.A1(new_n497_), .A2(new_n503_), .A3(new_n505_), .A4(new_n508_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n525_), .B(new_n527_), .C1(new_n533_), .C2(new_n526_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n450_), .B1(new_n521_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT106), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n511_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n537_), .A2(KEYINPUT27), .A3(new_n510_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT27), .B1(new_n510_), .B2(new_n515_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n450_), .A2(new_n536_), .A3(new_n524_), .A4(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n441_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n447_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n540_), .A2(new_n542_), .A3(new_n524_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT106), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n336_), .B1(new_n535_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT107), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n543_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n540_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT108), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n336_), .A2(new_n525_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(KEYINPUT107), .B(new_n336_), .C1(new_n535_), .C2(new_n546_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n549_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n269_), .B(KEYINPUT75), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT16), .B(G183gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT68), .B1(new_n561_), .B2(KEYINPUT17), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n557_), .B(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(new_n210_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(KEYINPUT17), .B2(new_n561_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT76), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n236_), .A2(new_n274_), .B1(new_n279_), .B2(new_n232_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(KEYINPUT35), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT34), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n235_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n234_), .B1(new_n224_), .B2(new_n231_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n274_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n279_), .A2(new_n232_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT34), .ZN(new_n581_));
  INV_X1    g380(.A(G232gat), .ZN(new_n582_));
  INV_X1    g381(.A(G233gat), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n575_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n575_), .B2(new_n581_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n572_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n574_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n580_), .A2(KEYINPUT34), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n584_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n575_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT35), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n588_), .A2(new_n593_), .A3(KEYINPUT72), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G134gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G162gat), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(KEYINPUT36), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT35), .ZN(new_n600_));
  INV_X1    g399(.A(new_n572_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT36), .B(new_n597_), .C1(new_n600_), .C2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n598_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n588_), .A2(new_n593_), .A3(KEYINPUT72), .A4(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n599_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT73), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(new_n607_), .A3(KEYINPUT37), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n569_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n260_), .A2(new_n294_), .A3(new_n556_), .A4(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n525_), .A3(new_n261_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n258_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n294_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n569_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n606_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n621_), .A2(new_n556_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n524_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(new_n625_), .ZN(G1324gat));
  OAI21_X1  g425(.A(G8gat), .B1(new_n624_), .B2(new_n540_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT39), .ZN(new_n628_));
  INV_X1    g427(.A(new_n540_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n615_), .A2(new_n262_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g431(.A(G15gat), .B1(new_n624_), .B2(new_n336_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT41), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n614_), .A2(G15gat), .A3(new_n336_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1326gat));
  OAI21_X1  g435(.A(G22gat), .B1(new_n624_), .B2(new_n550_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT42), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n614_), .A2(G22gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n550_), .B2(new_n639_), .ZN(G1327gat));
  AND3_X1   g439(.A1(new_n549_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(new_n623_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n622_), .A2(new_n620_), .A3(new_n619_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT114), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT114), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n646_), .A3(new_n643_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(G29gat), .B1(new_n648_), .B2(new_n525_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n606_), .A2(new_n607_), .A3(KEYINPUT37), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT37), .B1(new_n606_), .B2(new_n607_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT111), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT111), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n610_), .A2(new_n653_), .A3(new_n611_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n556_), .A2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n612_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(KEYINPUT43), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n656_), .A2(new_n658_), .B1(new_n556_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(KEYINPUT44), .A3(new_n643_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT112), .ZN(new_n665_));
  INV_X1    g464(.A(new_n643_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n661_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n660_), .A2(new_n556_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n657_), .B1(new_n556_), .B2(new_n655_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT112), .B(new_n643_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n668_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT113), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n667_), .A2(KEYINPUT113), .A3(new_n668_), .A4(new_n671_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n664_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(new_n525_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n649_), .B1(new_n677_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n645_), .A2(new_n679_), .A3(new_n629_), .A4(new_n647_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT45), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n663_), .A2(new_n629_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n683_), .B2(new_n679_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n681_), .B(KEYINPUT46), .C1(new_n683_), .C2(new_n679_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1329gat));
  NOR2_X1   g487(.A1(new_n336_), .A2(new_n271_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n664_), .B(new_n690_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n336_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G43gat), .B1(new_n648_), .B2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT47), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n676_), .A2(new_n689_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  INV_X1    g495(.A(new_n693_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n698_), .ZN(G1330gat));
  AOI21_X1  g498(.A(G50gat), .B1(new_n648_), .B2(new_n450_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n550_), .A2(new_n273_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n676_), .B2(new_n701_), .ZN(G1331gat));
  NAND2_X1  g501(.A1(new_n613_), .A2(new_n620_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n703_), .A2(new_n641_), .A3(new_n258_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n525_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n259_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n706_), .A2(new_n294_), .A3(new_n641_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n525_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n705_), .B1(new_n708_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g508(.A(G64gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n707_), .B2(new_n629_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT48), .Z(new_n712_));
  NOR2_X1   g511(.A1(new_n540_), .A2(G64gat), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT115), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n704_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1333gat));
  INV_X1    g515(.A(G71gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n707_), .B2(new_n692_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT49), .Z(new_n719_));
  NAND3_X1  g518(.A1(new_n704_), .A2(new_n717_), .A3(new_n692_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1334gat));
  NOR2_X1   g520(.A1(new_n550_), .A2(G78gat), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT116), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n704_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n707_), .A2(new_n450_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G78gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G78gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT117), .Z(G1335gat));
  NOR2_X1   g529(.A1(new_n622_), .A2(new_n294_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n642_), .A2(new_n259_), .A3(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT118), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n525_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n662_), .A2(new_n619_), .A3(new_n731_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(new_n524_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(G85gat), .B2(new_n736_), .ZN(G1336gat));
  AOI21_X1  g536(.A(G92gat), .B1(new_n733_), .B2(new_n629_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n735_), .A2(new_n540_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(G92gat), .B2(new_n739_), .ZN(G1337gat));
  NAND3_X1  g539(.A1(new_n733_), .A2(new_n227_), .A3(new_n692_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G99gat), .B1(new_n735_), .B2(new_n336_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n228_), .A3(new_n450_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n662_), .A2(new_n619_), .A3(new_n450_), .A4(new_n731_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n746_), .B2(G106gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n745_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g551(.A(KEYINPUT57), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n242_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n244_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n241_), .A2(KEYINPUT55), .A3(new_n242_), .A4(new_n243_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n253_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n247_), .A2(new_n254_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n294_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n756_), .A2(new_n757_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n253_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n758_), .A2(KEYINPUT56), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n283_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n281_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n276_), .A2(new_n283_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n291_), .A3(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n293_), .A2(new_n771_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n761_), .A2(new_n767_), .B1(new_n255_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n753_), .B1(new_n773_), .B2(new_n606_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n761_), .A2(new_n767_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n255_), .A2(new_n772_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT57), .B(new_n623_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n778_));
  INV_X1    g577(.A(new_n760_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n772_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n780_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n772_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n612_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n774_), .B(new_n777_), .C1(new_n785_), .C2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n569_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT54), .B1(new_n703_), .B2(new_n619_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n613_), .A2(new_n791_), .A3(new_n620_), .A4(new_n258_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(new_n525_), .A3(new_n552_), .A4(new_n692_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G113gat), .B1(new_n796_), .B2(new_n294_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(KEYINPUT121), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n795_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(KEYINPUT121), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n795_), .B2(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n800_), .A2(new_n802_), .A3(new_n620_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n797_), .B1(new_n803_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g603(.A(new_n333_), .B1(new_n258_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n796_), .B(new_n805_), .C1(KEYINPUT60), .C2(new_n333_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n800_), .A2(new_n802_), .A3(new_n260_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n333_), .ZN(G1341gat));
  AOI21_X1  g607(.A(G127gat), .B1(new_n796_), .B2(new_n622_), .ZN(new_n809_));
  INV_X1    g608(.A(G127gat), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n800_), .A2(new_n802_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n811_), .B2(new_n622_), .ZN(G1342gat));
  AOI21_X1  g611(.A(G134gat), .B1(new_n796_), .B2(new_n606_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n800_), .A2(new_n802_), .A3(new_n659_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(G134gat), .ZN(G1343gat));
  AOI22_X1  g614(.A1(new_n569_), .A2(new_n788_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n816_), .A2(new_n524_), .A3(new_n629_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n692_), .A2(new_n550_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n620_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(new_n351_), .ZN(G1344gat));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n260_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(new_n352_), .ZN(G1345gat));
  AND2_X1   g622(.A1(new_n817_), .A2(new_n818_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n622_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT61), .B(G155gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(G1346gat));
  AOI21_X1  g626(.A(G162gat), .B1(new_n824_), .B2(new_n606_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n655_), .A2(G162gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n824_), .B2(new_n829_), .ZN(G1347gat));
  NOR2_X1   g629(.A1(new_n816_), .A2(new_n450_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n553_), .A2(new_n629_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n620_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n318_), .A3(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n833_), .B(KEYINPUT122), .Z(new_n835_));
  AOI21_X1  g634(.A(new_n289_), .B1(new_n831_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n837_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n834_), .B1(new_n838_), .B2(new_n839_), .ZN(G1348gat));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n816_), .B2(new_n450_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n794_), .A2(KEYINPUT123), .A3(new_n550_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n832_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n842_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n845_), .A2(KEYINPUT124), .A3(G176gat), .A4(new_n259_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n831_), .A2(new_n844_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n252_), .B1(new_n847_), .B2(new_n258_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n842_), .A2(new_n843_), .A3(G176gat), .A4(new_n844_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n260_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n846_), .A2(new_n848_), .A3(new_n851_), .ZN(G1349gat));
  AOI21_X1  g651(.A(G183gat), .B1(new_n845_), .B2(new_n622_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n847_), .A2(new_n569_), .A3(new_n298_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n847_), .B2(new_n659_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n606_), .A2(new_n299_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n847_), .B2(new_n857_), .ZN(G1351gat));
  NOR2_X1   g657(.A1(new_n550_), .A2(new_n525_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n692_), .A2(new_n540_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n794_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n620_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n407_), .ZN(G1352gat));
  AND3_X1   g662(.A1(new_n794_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n259_), .A3(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT126), .Z(new_n868_));
  XNOR2_X1  g667(.A(new_n866_), .B(new_n868_), .ZN(G1353gat));
  NAND2_X1  g668(.A1(new_n864_), .A2(new_n622_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  AND2_X1   g670(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n870_), .B2(new_n871_), .ZN(G1354gat));
  INV_X1    g673(.A(G218gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n864_), .A2(new_n875_), .A3(new_n606_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G218gat), .B1(new_n861_), .B2(new_n659_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


