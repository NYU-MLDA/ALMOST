//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n973_, new_n974_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n991_, new_n992_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n999_, new_n1000_;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203_));
  INV_X1    g002(.A(G85gat), .ZN(new_n204_));
  INV_X1    g003(.A(G92gat), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT9), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  AOI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(KEYINPUT9), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT10), .B(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(new_n211_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT64), .B(KEYINPUT6), .Z(new_n217_));
  INV_X1    g016(.A(new_n215_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n208_), .A2(new_n212_), .A3(new_n216_), .A4(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  OAI22_X1  g020(.A1(new_n221_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  OR4_X1    g021(.A1(new_n221_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n219_), .A2(new_n216_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n224_), .A2(new_n207_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(new_n224_), .B2(new_n207_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n220_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT69), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n230_), .B(new_n220_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G29gat), .B(G36gat), .Z(new_n232_));
  XOR2_X1   g031(.A(G43gat), .B(G50gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT15), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n229_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G232gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT34), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT35), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n220_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n227_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n224_), .A2(new_n207_), .A3(new_n225_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n246_), .A2(new_n234_), .B1(new_n240_), .B2(new_n239_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n236_), .A2(new_n242_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n242_), .B1(new_n236_), .B2(new_n247_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n203_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n236_), .A2(new_n247_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n241_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n236_), .A2(new_n247_), .A3(new_n242_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT75), .A3(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G190gat), .B(G218gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT71), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G134gat), .B(G162gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT36), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(new_n254_), .A3(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n248_), .A2(new_n249_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT36), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT72), .B1(new_n261_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n266_));
  NOR4_X1   g065(.A1(new_n248_), .A2(new_n249_), .A3(new_n266_), .A4(new_n263_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n260_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n261_), .A2(KEYINPUT72), .A3(new_n264_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n252_), .A2(new_n264_), .A3(new_n253_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n266_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n259_), .B(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(KEYINPUT74), .B(new_n276_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n276_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n274_), .A2(KEYINPUT37), .A3(new_n277_), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n270_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G127gat), .B(G155gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G183gat), .B(G211gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT17), .ZN(new_n288_));
  INV_X1    g087(.A(G231gat), .ZN(new_n289_));
  INV_X1    g088(.A(G233gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT76), .B(G8gat), .ZN(new_n292_));
  INV_X1    g091(.A(G1gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT14), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT77), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n298_), .A3(new_n295_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n291_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(new_n299_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n300_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n291_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n301_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G71gat), .B(G78gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G57gat), .B(G64gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT67), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n314_), .B2(KEYINPUT11), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n313_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT11), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n317_), .A2(KEYINPUT68), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n314_), .B2(KEYINPUT11), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n315_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT68), .B1(new_n317_), .B2(new_n318_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n311_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n314_), .A2(new_n320_), .A3(KEYINPUT11), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n310_), .A2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n304_), .A2(new_n309_), .A3(new_n326_), .A4(new_n322_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n288_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n287_), .A2(KEYINPUT17), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT79), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n328_), .A2(new_n329_), .A3(new_n334_), .A4(new_n331_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n330_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n202_), .B1(new_n282_), .B2(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n280_), .A2(new_n277_), .A3(KEYINPUT37), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n274_), .A2(new_n339_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT80), .A3(new_n336_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT13), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n327_), .A2(new_n228_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n327_), .A2(new_n228_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT12), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G230gat), .A2(G233gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n229_), .A2(KEYINPUT12), .A3(new_n327_), .A4(new_n231_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n345_), .ZN(new_n352_));
  OAI211_X1 g151(.A(G230gat), .B(G233gat), .C1(new_n352_), .C2(new_n346_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G120gat), .B(G148gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT5), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G176gat), .B(G204gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT70), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n351_), .A2(new_n353_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n344_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n351_), .A2(new_n353_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT13), .A3(new_n359_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n342_), .A2(new_n343_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n338_), .A2(new_n341_), .A3(new_n367_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT81), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  INV_X1    g172(.A(G197gat), .ZN(new_n374_));
  INV_X1    g173(.A(G204gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G197gat), .A2(G204gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(KEYINPUT21), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G211gat), .B(G218gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT91), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n377_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G197gat), .A2(G204gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT21), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT91), .ZN(new_n385_));
  XOR2_X1   g184(.A(G211gat), .B(G218gat), .Z(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n378_), .A2(new_n379_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n380_), .A2(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G183gat), .ZN(new_n391_));
  INV_X1    g190(.A(G190gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT23), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G183gat), .A3(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G169gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G169gat), .A2(G176gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT24), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT84), .B1(new_n392_), .B2(KEYINPUT26), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT26), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(G190gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n391_), .A2(KEYINPUT25), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT25), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G183gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n392_), .A2(KEYINPUT26), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(KEYINPUT85), .B(new_n405_), .C1(new_n410_), .C2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n395_), .A2(KEYINPUT86), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n395_), .A2(KEYINPUT86), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n393_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n403_), .A2(KEYINPUT24), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT25), .B(G183gat), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n422_), .A2(new_n414_), .A3(new_n406_), .A4(new_n409_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT85), .B1(new_n423_), .B2(new_n405_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n390_), .B(new_n402_), .C1(new_n421_), .C2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT20), .ZN(new_n427_));
  INV_X1    g226(.A(new_n390_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n420_), .A2(new_n396_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G190gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n422_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n405_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT95), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(KEYINPUT95), .A3(new_n405_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n429_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n401_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n419_), .B2(new_n398_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n428_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n427_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n426_), .B1(new_n425_), .B2(KEYINPUT20), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n373_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT18), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n434_), .A2(new_n435_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n429_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n438_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n390_), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n402_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n428_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n373_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT20), .A4(new_n455_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n442_), .A2(new_n447_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n447_), .B1(new_n442_), .B2(new_n456_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n371_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n440_), .A2(new_n373_), .A3(new_n441_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n450_), .A2(KEYINPUT101), .A3(new_n451_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT101), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n390_), .A3(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n453_), .B2(new_n428_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n455_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n446_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n442_), .A2(new_n447_), .A3(new_n456_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT27), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n459_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G22gat), .B(G50gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT28), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G141gat), .A2(G148gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(KEYINPUT3), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT3), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(KEYINPUT89), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT2), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT2), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G141gat), .A3(G148gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(G141gat), .A2(G148gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(KEYINPUT90), .A3(KEYINPUT3), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n480_), .A2(new_n485_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n492_));
  INV_X1    g291(.A(G155gat), .ZN(new_n493_));
  INV_X1    g292(.A(G162gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n495_), .A2(new_n496_), .B1(G155gat), .B2(G162gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G155gat), .A2(G162gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT1), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n489_), .A2(new_n481_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n491_), .A2(new_n497_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT29), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n474_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n498_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n478_), .A2(KEYINPUT89), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n476_), .A2(KEYINPUT3), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n511_), .A2(new_n475_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n486_), .B(KEYINPUT90), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n508_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n503_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n515_));
  NOR4_X1   g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n473_), .B1(new_n507_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT89), .B(KEYINPUT3), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n485_), .B1(new_n519_), .B2(new_n489_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n490_), .A2(new_n488_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n497_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n502_), .A2(new_n504_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n506_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT28), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n505_), .A2(new_n474_), .A3(new_n506_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n472_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n517_), .A2(new_n518_), .A3(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT29), .B1(new_n514_), .B2(new_n515_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G228gat), .A2(G233gat), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n428_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n428_), .B2(new_n529_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G78gat), .B(G106gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n517_), .A2(new_n527_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT93), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT92), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(new_n540_), .A3(KEYINPUT93), .ZN(new_n541_));
  INV_X1    g340(.A(new_n535_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n528_), .A2(new_n542_), .A3(new_n533_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n536_), .A2(new_n539_), .A3(new_n541_), .A4(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n528_), .A2(new_n542_), .A3(new_n533_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n540_), .B1(new_n537_), .B2(KEYINPUT93), .ZN(new_n547_));
  AOI211_X1 g346(.A(KEYINPUT92), .B(new_n518_), .C1(new_n517_), .C2(new_n527_), .ZN(new_n548_));
  OAI22_X1  g347(.A1(new_n545_), .A2(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n544_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G85gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT98), .Z(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n293_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n551_), .B(KEYINPUT98), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G1gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n557_));
  INV_X1    g356(.A(G29gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n553_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G127gat), .B(G134gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G113gat), .B(G120gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n564_), .B(new_n565_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n522_), .A2(new_n568_), .A3(new_n523_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n569_), .A3(KEYINPUT4), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G225gat), .A2(G233gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT4), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n566_), .B(new_n574_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .A4(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n567_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n573_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n571_), .B1(new_n580_), .B2(new_n570_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n563_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n567_), .A2(KEYINPUT4), .A3(new_n569_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT96), .B1(new_n583_), .B2(new_n579_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n563_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n577_), .A4(new_n576_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G71gat), .B(G99gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(G43gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n453_), .B(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G227gat), .A2(G233gat), .ZN(new_n595_));
  INV_X1    g394(.A(G15gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT30), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(new_n566_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n593_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n594_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n594_), .B2(new_n600_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n588_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n471_), .A2(new_n550_), .A3(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n550_), .A2(new_n459_), .A3(new_n588_), .A4(new_n470_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n457_), .A2(new_n458_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n578_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n585_), .A4(new_n584_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n586_), .A2(KEYINPUT33), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n567_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n563_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT99), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n570_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n612_), .B2(KEYINPUT99), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n609_), .A2(new_n610_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n456_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n425_), .A2(KEYINPUT20), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT94), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n439_), .A3(new_n427_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n617_), .B1(new_n620_), .B2(new_n373_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n447_), .A2(KEYINPUT32), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n621_), .A2(new_n622_), .B1(new_n582_), .B2(new_n586_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n606_), .A2(new_n616_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n605_), .B1(new_n626_), .B2(new_n550_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n601_), .A2(new_n602_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n604_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n234_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT82), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n307_), .A2(new_n301_), .A3(new_n234_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(KEYINPUT82), .B(new_n630_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n235_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n635_), .A3(new_n633_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT83), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G169gat), .B(G197gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n638_), .A2(new_n640_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n629_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n368_), .A2(new_n370_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n368_), .A2(KEYINPUT102), .A3(new_n370_), .A4(new_n649_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n588_), .A2(G1gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(KEYINPUT38), .A3(new_n655_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n268_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n629_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n362_), .A2(new_n366_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n648_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n336_), .A3(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n588_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n658_), .A2(new_n659_), .A3(new_n665_), .ZN(G1324gat));
  NAND4_X1  g465(.A1(new_n652_), .A2(new_n292_), .A3(new_n471_), .A4(new_n653_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n442_), .A2(new_n456_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n446_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n469_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n371_), .B1(new_n621_), .B2(new_n447_), .ZN(new_n672_));
  AOI22_X1  g471(.A1(new_n671_), .A2(new_n371_), .B1(new_n672_), .B2(new_n468_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G8gat), .B1(new_n664_), .B2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n668_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n667_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n667_), .A2(new_n678_), .A3(KEYINPUT40), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1325gat));
  INV_X1    g482(.A(new_n628_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n654_), .A2(new_n596_), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G15gat), .B1(new_n664_), .B2(new_n628_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(KEYINPUT104), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(KEYINPUT104), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(KEYINPUT41), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(KEYINPUT41), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n685_), .B1(new_n690_), .B2(new_n691_), .ZN(G1326gat));
  INV_X1    g491(.A(new_n550_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(G22gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n654_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G22gat), .B1(new_n664_), .B2(new_n693_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT42), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1327gat));
  NOR3_X1   g498(.A1(new_n662_), .A2(new_n336_), .A3(new_n268_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n649_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n558_), .A3(new_n587_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n629_), .B2(new_n340_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n625_), .B(new_n587_), .C1(new_n669_), .C2(new_n624_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n609_), .A2(new_n610_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n613_), .A2(new_n615_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n709_), .B2(new_n671_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n693_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n684_), .B1(new_n711_), .B2(new_n605_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n705_), .B(new_n282_), .C1(new_n712_), .C2(new_n604_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n704_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n663_), .A2(new_n337_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  AOI211_X1 g517(.A(new_n718_), .B(new_n715_), .C1(new_n704_), .C2(new_n713_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n587_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n721_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT106), .B1(new_n721_), .B2(G29gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n703_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n725_), .A2(KEYINPUT108), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n673_), .A2(G36gat), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n701_), .A2(KEYINPUT45), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT45), .B1(new_n701_), .B2(new_n727_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n728_), .A2(new_n729_), .B1(KEYINPUT108), .B2(new_n725_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n604_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n587_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n732_));
  AOI22_X1  g531(.A1(new_n710_), .A2(new_n693_), .B1(new_n673_), .B2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n733_), .B2(new_n684_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n705_), .B1(new_n734_), .B2(new_n282_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n629_), .A2(KEYINPUT43), .A3(new_n340_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n716_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n718_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n714_), .A2(KEYINPUT44), .A3(new_n716_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n738_), .A2(KEYINPUT107), .A3(new_n471_), .A4(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G36gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT107), .B1(new_n720_), .B2(new_n471_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n726_), .B(new_n730_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n738_), .A2(new_n471_), .A3(new_n739_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(G36gat), .A3(new_n740_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n726_), .B1(new_n748_), .B2(new_n730_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n744_), .A2(new_n749_), .ZN(G1329gat));
  NOR3_X1   g549(.A1(new_n717_), .A2(new_n719_), .A3(new_n628_), .ZN(new_n751_));
  INV_X1    g550(.A(G43gat), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n684_), .A2(new_n752_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n701_), .A2(new_n755_), .ZN(new_n756_));
  OR3_X1    g555(.A1(new_n753_), .A2(new_n754_), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n753_), .B2(new_n756_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1330gat));
  AOI21_X1  g558(.A(G50gat), .B1(new_n702_), .B2(new_n550_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n550_), .A2(G50gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n720_), .B2(new_n761_), .ZN(G1331gat));
  INV_X1    g561(.A(new_n648_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n629_), .A2(new_n367_), .A3(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n342_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n587_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n661_), .A2(new_n662_), .A3(new_n336_), .A4(new_n648_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G57gat), .B1(new_n768_), .B2(new_n588_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1332gat));
  OAI21_X1  g569(.A(G64gat), .B1(new_n768_), .B2(new_n673_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT48), .ZN(new_n772_));
  INV_X1    g571(.A(G64gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n773_), .A3(new_n471_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n768_), .B2(new_n628_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT109), .B(KEYINPUT49), .Z(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(G71gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n779_), .A3(new_n684_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1334gat));
  OAI21_X1  g580(.A(G78gat), .B1(new_n768_), .B2(new_n693_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT50), .ZN(new_n783_));
  INV_X1    g582(.A(G78gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n765_), .A2(new_n784_), .A3(new_n550_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n268_), .A2(new_n336_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n764_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(G85gat), .B1(new_n789_), .B2(new_n587_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n367_), .A2(new_n763_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n714_), .A2(new_n337_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n587_), .A2(G85gat), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT110), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n790_), .B1(new_n793_), .B2(new_n795_), .ZN(G1336gat));
  OAI21_X1  g595(.A(G92gat), .B1(new_n792_), .B2(new_n673_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n789_), .A2(new_n205_), .A3(new_n471_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n792_), .B2(new_n628_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n684_), .A2(new_n210_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n788_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g602(.A1(new_n789_), .A2(new_n211_), .A3(new_n550_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n793_), .A2(new_n550_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(G106gat), .ZN(new_n807_));
  AOI211_X1 g606(.A(KEYINPUT52), .B(new_n211_), .C1(new_n793_), .C2(new_n550_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n804_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  NAND2_X1  g612(.A1(new_n648_), .A2(new_n336_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n648_), .A2(new_n336_), .A3(KEYINPUT111), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n367_), .A2(new_n818_), .A3(new_n270_), .A4(new_n281_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT112), .B1(new_n819_), .B2(KEYINPUT54), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n648_), .A2(new_n336_), .A3(KEYINPUT111), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT111), .B1(new_n648_), .B2(new_n336_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n366_), .B(new_n362_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n282_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n282_), .B2(new_n823_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT113), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n819_), .A2(new_n830_), .A3(KEYINPUT54), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n820_), .A2(new_n827_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n363_), .A2(new_n357_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n633_), .A2(new_n636_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n644_), .B1(new_n834_), .B2(new_n639_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n634_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n645_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n645_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT114), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n833_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n349_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n351_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n348_), .A2(KEYINPUT55), .A3(new_n349_), .A4(new_n350_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n357_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  INV_X1    g648(.A(new_n357_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n849_), .B(new_n850_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n842_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI221_X1 g653(.A(new_n842_), .B1(KEYINPUT115), .B2(KEYINPUT58), .C1(new_n848_), .C2(new_n851_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n282_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT116), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n854_), .A2(new_n855_), .A3(new_n858_), .A4(new_n282_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n833_), .A2(new_n648_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n847_), .A2(new_n357_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n849_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n357_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n841_), .A2(new_n839_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n360_), .A2(new_n361_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n268_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n860_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n868_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(KEYINPUT57), .A3(new_n268_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n857_), .A2(new_n859_), .A3(new_n871_), .A4(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n832_), .B1(new_n876_), .B2(new_n337_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n471_), .A2(new_n550_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n587_), .A3(new_n684_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n877_), .A2(new_n648_), .A3(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT117), .B1(new_n880_), .B2(G113gat), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882_));
  INV_X1    g681(.A(G113gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n876_), .A2(new_n337_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n832_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n879_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n882_), .B(new_n883_), .C1(new_n888_), .C2(new_n648_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n871_), .A2(new_n856_), .A3(new_n875_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n827_), .A2(new_n820_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n829_), .A2(new_n831_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n890_), .A2(new_n337_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n887_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n888_), .B2(KEYINPUT59), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n648_), .A2(new_n883_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT118), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n881_), .A2(new_n889_), .B1(new_n897_), .B2(new_n899_), .ZN(G1340gat));
  OR2_X1    g699(.A1(new_n893_), .A2(new_n895_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n877_), .A2(new_n879_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n662_), .B(new_n901_), .C1(new_n902_), .C2(new_n894_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G120gat), .ZN(new_n904_));
  INV_X1    g703(.A(G120gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n367_), .B2(KEYINPUT60), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n902_), .B(new_n906_), .C1(KEYINPUT60), .C2(new_n905_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(G1341gat));
  AOI21_X1  g707(.A(G127gat), .B1(new_n902_), .B2(new_n336_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n336_), .A2(G127gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT119), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n897_), .B2(new_n911_), .ZN(G1342gat));
  AOI21_X1  g711(.A(G134gat), .B1(new_n902_), .B2(new_n660_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n282_), .A2(G134gat), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT120), .Z(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n897_), .B2(new_n915_), .ZN(G1343gat));
  NOR4_X1   g715(.A1(new_n471_), .A2(new_n693_), .A3(new_n684_), .A4(new_n588_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n763_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n662_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g722(.A1(new_n886_), .A2(new_n336_), .A3(new_n917_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT121), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n919_), .A2(new_n926_), .A3(new_n336_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT61), .B(G155gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n925_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n928_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n926_), .B1(new_n919_), .B2(new_n336_), .ZN(new_n931_));
  NOR4_X1   g730(.A1(new_n877_), .A2(KEYINPUT121), .A3(new_n337_), .A4(new_n918_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n929_), .A2(new_n933_), .ZN(G1346gat));
  INV_X1    g733(.A(new_n919_), .ZN(new_n935_));
  OAI21_X1  g734(.A(G162gat), .B1(new_n935_), .B2(new_n340_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n919_), .A2(new_n494_), .A3(new_n660_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n673_), .A2(new_n603_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n693_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n893_), .A2(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n942_));
  AND2_X1   g741(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n941_), .B(new_n763_), .C1(new_n942_), .C2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n939_), .A2(new_n763_), .ZN(new_n946_));
  XOR2_X1   g745(.A(new_n946_), .B(KEYINPUT122), .Z(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n550_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n945_), .B1(new_n893_), .B2(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(KEYINPUT57), .B1(new_n874_), .B2(new_n268_), .ZN(new_n951_));
  AOI211_X1 g750(.A(new_n870_), .B(new_n660_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n336_), .B1(new_n953_), .B2(new_n856_), .ZN(new_n954_));
  OAI211_X1 g753(.A(KEYINPUT123), .B(new_n948_), .C1(new_n954_), .C2(new_n832_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n950_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957_));
  OAI21_X1  g756(.A(G169gat), .B1(new_n957_), .B2(KEYINPUT124), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  AOI22_X1  g758(.A1(new_n956_), .A2(new_n959_), .B1(KEYINPUT124), .B2(new_n957_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n957_), .A2(KEYINPUT124), .ZN(new_n961_));
  AOI211_X1 g760(.A(new_n961_), .B(new_n958_), .C1(new_n950_), .C2(new_n955_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n944_), .B1(new_n960_), .B2(new_n962_), .ZN(G1348gat));
  NAND3_X1  g762(.A1(new_n886_), .A2(KEYINPUT125), .A3(new_n693_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n965_), .B1(new_n877_), .B2(new_n550_), .ZN(new_n966_));
  INV_X1    g765(.A(G176gat), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n367_), .A2(new_n967_), .ZN(new_n968_));
  NAND4_X1  g767(.A1(new_n964_), .A2(new_n966_), .A3(new_n939_), .A4(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n941_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n967_), .B1(new_n970_), .B2(new_n367_), .ZN(new_n971_));
  AND2_X1   g770(.A1(new_n969_), .A2(new_n971_), .ZN(G1349gat));
  NOR3_X1   g771(.A1(new_n970_), .A2(new_n337_), .A3(new_n422_), .ZN(new_n973_));
  NAND4_X1  g772(.A1(new_n964_), .A2(new_n966_), .A3(new_n336_), .A4(new_n939_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n974_), .B2(new_n391_), .ZN(G1350gat));
  NAND2_X1  g774(.A1(new_n660_), .A2(new_n430_), .ZN(new_n976_));
  XOR2_X1   g775(.A(new_n976_), .B(KEYINPUT126), .Z(new_n977_));
  NAND2_X1  g776(.A1(new_n941_), .A2(new_n977_), .ZN(new_n978_));
  NOR3_X1   g777(.A1(new_n893_), .A2(new_n340_), .A3(new_n940_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n392_), .B2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n980_), .A2(KEYINPUT127), .ZN(new_n981_));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982_));
  OAI211_X1 g781(.A(new_n978_), .B(new_n982_), .C1(new_n392_), .C2(new_n979_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n981_), .A2(new_n983_), .ZN(G1351gat));
  AND3_X1   g783(.A1(new_n471_), .A2(new_n732_), .A3(new_n628_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n886_), .A2(new_n985_), .ZN(new_n986_));
  INV_X1    g785(.A(new_n986_), .ZN(new_n987_));
  AOI21_X1  g786(.A(G197gat), .B1(new_n987_), .B2(new_n763_), .ZN(new_n988_));
  NOR3_X1   g787(.A1(new_n986_), .A2(new_n374_), .A3(new_n648_), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n988_), .A2(new_n989_), .ZN(G1352gat));
  NAND3_X1  g789(.A1(new_n987_), .A2(new_n375_), .A3(new_n662_), .ZN(new_n991_));
  OAI21_X1  g790(.A(G204gat), .B1(new_n986_), .B2(new_n367_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n991_), .A2(new_n992_), .ZN(G1353gat));
  XNOR2_X1  g792(.A(KEYINPUT63), .B(G211gat), .ZN(new_n994_));
  NOR3_X1   g793(.A1(new_n986_), .A2(new_n337_), .A3(new_n994_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n987_), .A2(new_n336_), .ZN(new_n996_));
  NOR2_X1   g795(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n995_), .B1(new_n996_), .B2(new_n997_), .ZN(G1354gat));
  OR3_X1    g797(.A1(new_n986_), .A2(G218gat), .A3(new_n268_), .ZN(new_n999_));
  OAI21_X1  g798(.A(G218gat), .B1(new_n986_), .B2(new_n340_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n999_), .A2(new_n1000_), .ZN(G1355gat));
endmodule


