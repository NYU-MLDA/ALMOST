//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n969_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1009_, new_n1010_, new_n1011_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1031_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1042_,
    new_n1043_, new_n1044_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT96), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT93), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT25), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n212_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(KEYINPUT25), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(G183gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT93), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT94), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n222_), .A2(new_n223_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n223_), .B1(new_n222_), .B2(new_n228_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT79), .ZN(new_n233_));
  OR3_X1    g032(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n234_));
  INV_X1    g033(.A(G190gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT23), .B1(new_n215_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n232_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT79), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n233_), .B(new_n234_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n229_), .A2(new_n230_), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G169gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n211_), .B1(new_n240_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n222_), .A2(new_n228_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n239_), .B1(new_n248_), .B2(KEYINPUT94), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n222_), .A2(new_n223_), .A3(new_n228_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n246_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT96), .ZN(new_n252_));
  INV_X1    g051(.A(G218gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G211gat), .ZN(new_n254_));
  INV_X1    g053(.A(G211gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G218gat), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT90), .ZN(new_n262_));
  INV_X1    g061(.A(G197gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(G204gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT21), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(KEYINPUT90), .B2(new_n259_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(G204gat), .ZN(new_n267_));
  INV_X1    g066(.A(G204gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(G197gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n257_), .B1(new_n270_), .B2(KEYINPUT21), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n261_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n254_), .A2(new_n256_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n274_));
  OAI211_X1 g073(.A(KEYINPUT21), .B(new_n264_), .C1(new_n270_), .C2(new_n262_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT91), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n260_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n247_), .A2(new_n252_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT20), .ZN(new_n279_));
  INV_X1    g078(.A(new_n260_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT91), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT91), .B1(new_n274_), .B2(new_n275_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n237_), .A2(new_n228_), .A3(new_n234_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT25), .B(G183gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(new_n218_), .A3(KEYINPUT78), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT78), .B1(new_n285_), .B2(new_n218_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n284_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n233_), .B(new_n241_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n244_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n279_), .B1(new_n283_), .B2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n210_), .B1(new_n278_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n248_), .A2(KEYINPUT94), .ZN(new_n295_));
  INV_X1    g094(.A(new_n239_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n250_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n277_), .B1(new_n297_), .B2(new_n245_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT20), .B1(new_n283_), .B2(new_n292_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n209_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n207_), .B1(new_n294_), .B2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n209_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(new_n277_), .A3(new_n245_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n293_), .A2(new_n303_), .A3(new_n210_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n206_), .A3(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n305_), .A2(KEYINPUT27), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n283_), .B1(new_n240_), .B2(new_n246_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n285_), .A2(new_n218_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n286_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n311_), .A2(new_n284_), .B1(new_n290_), .B2(new_n244_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n279_), .B1(new_n277_), .B2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n210_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n297_), .A2(new_n277_), .A3(new_n245_), .ZN(new_n315_));
  OAI211_X1 g114(.A(KEYINPUT20), .B(new_n210_), .C1(new_n277_), .C2(new_n312_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n207_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n305_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT27), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n301_), .A2(new_n306_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT86), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n330_), .B(new_n331_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n337_), .A2(KEYINPUT86), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT85), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT85), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT3), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(G141gat), .B2(G148gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n344_), .A2(G141gat), .A3(G148gat), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n341_), .B(new_n343_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n329_), .B1(new_n339_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n335_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n325_), .A2(KEYINPUT1), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n325_), .B1(new_n327_), .B2(KEYINPUT1), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT83), .B(new_n325_), .C1(new_n327_), .C2(KEYINPUT1), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n353_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n324_), .B1(new_n349_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n341_), .A2(new_n343_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n347_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(new_n345_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n337_), .A2(KEYINPUT86), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n332_), .A2(new_n333_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n330_), .A4(new_n331_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n328_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n355_), .A2(new_n356_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n354_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n358_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n352_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n371_), .A3(KEYINPUT87), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n360_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n323_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G22gat), .B(G50gat), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n373_), .A2(new_n374_), .A3(new_n323_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI211_X1 g179(.A(KEYINPUT29), .B(new_n322_), .C1(new_n360_), .C2(new_n372_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n377_), .B1(new_n375_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n360_), .A2(new_n372_), .A3(KEYINPUT29), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT89), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n360_), .A2(new_n372_), .A3(new_n386_), .A4(KEYINPUT29), .ZN(new_n387_));
  AND2_X1   g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n277_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n277_), .B2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G78gat), .B(G106gat), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n390_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n383_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n384_), .A2(KEYINPUT89), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n387_), .A2(new_n389_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n393_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n394_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n390_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n402_), .A2(new_n382_), .A3(new_n380_), .A4(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n321_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n292_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n312_), .A2(KEYINPUT30), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G71gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G99gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n410_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(G127gat), .B(G134gat), .Z(new_n421_));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G127gat), .B(G134gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT81), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n425_), .A3(new_n420_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n419_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n428_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n431_), .A2(new_n426_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT80), .B(G43gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT31), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n436_), .A3(new_n433_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n360_), .A2(new_n372_), .A3(new_n432_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n429_), .A2(new_n371_), .A3(new_n367_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n449_), .B2(new_n442_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G85gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT0), .B(G57gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n443_), .A2(new_n444_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT4), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n443_), .A2(new_n446_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n442_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n445_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n454_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n406_), .A2(new_n440_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT97), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n398_), .A2(new_n404_), .A3(new_n455_), .A4(new_n463_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n302_), .A2(new_n206_), .A3(new_n304_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n206_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n320_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n277_), .B1(new_n251_), .B2(KEYINPUT96), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n240_), .A2(new_n211_), .A3(new_n246_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n293_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n209_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n300_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n206_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n305_), .A2(KEYINPUT27), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n470_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n466_), .B1(new_n467_), .B2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n398_), .A2(new_n404_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n459_), .A2(new_n454_), .A3(new_n460_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n454_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n480_), .A2(new_n321_), .A3(KEYINPUT97), .A4(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT33), .B1(new_n461_), .B2(new_n462_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n441_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n443_), .A2(new_n444_), .A3(new_n442_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n487_), .A2(new_n454_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(new_n305_), .A3(new_n318_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n482_), .A2(KEYINPUT33), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n302_), .A2(new_n304_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n474_), .A2(new_n475_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(new_n494_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n491_), .A2(new_n492_), .B1(new_n497_), .B2(new_n464_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n479_), .B(new_n484_), .C1(new_n498_), .C2(new_n480_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n438_), .A2(new_n439_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT82), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n465_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G169gat), .B(G197gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G1gat), .B(G8gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT14), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT74), .B(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n512_), .B2(G8gat), .ZN(new_n513_));
  OR2_X1    g312(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G22gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(G22gat), .A3(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n509_), .B1(new_n513_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n523_), .A2(new_n519_), .A3(new_n518_), .A4(new_n508_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT71), .ZN(new_n525_));
  INV_X1    g324(.A(G29gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(G36gat), .ZN(new_n527_));
  INV_X1    g326(.A(G36gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(G29gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n525_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(G29gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(G36gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT71), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n530_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT71), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT71), .B1(new_n531_), .B2(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n521_), .A2(new_n524_), .A3(new_n535_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n521_), .A2(new_n524_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n507_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(KEYINPUT77), .A3(new_n540_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n539_), .A2(new_n535_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT15), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(new_n524_), .A3(new_n521_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(new_n546_), .A3(new_n544_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n506_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n548_), .A2(new_n552_), .A3(new_n506_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n503_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561_));
  INV_X1    g360(.A(G99gat), .ZN(new_n562_));
  INV_X1    g361(.A(G106gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT6), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(G99gat), .B2(G106gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(KEYINPUT6), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n560_), .B(new_n564_), .C1(new_n566_), .C2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT64), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(KEYINPUT8), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(KEYINPUT8), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n569_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n572_), .B1(new_n569_), .B2(new_n577_), .ZN(new_n579_));
  OR2_X1    g378(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n563_), .A3(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n573_), .A2(KEYINPUT9), .A3(new_n575_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n567_), .A2(KEYINPUT6), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n565_), .A2(G99gat), .A3(G106gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n575_), .A2(KEYINPUT9), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n582_), .A2(new_n583_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n578_), .A2(new_n579_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT66), .ZN(new_n591_));
  INV_X1    g390(.A(G71gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT65), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT65), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(G71gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(G78gat), .ZN(new_n597_));
  INV_X1    g396(.A(G78gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(G64gat), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(G57gat), .ZN(new_n601_));
  INV_X1    g400(.A(G57gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(G64gat), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n601_), .A2(new_n603_), .A3(KEYINPUT11), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT11), .B1(new_n601_), .B2(new_n603_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n597_), .B(new_n599_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n603_), .A3(KEYINPUT11), .ZN(new_n607_));
  INV_X1    g406(.A(new_n599_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n598_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n590_), .A2(new_n591_), .A3(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n584_), .A2(new_n585_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n564_), .A2(new_n560_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n577_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n571_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n569_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n588_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT66), .B1(new_n619_), .B2(new_n611_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n613_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n590_), .A2(new_n612_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n559_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT12), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(new_n590_), .B2(new_n612_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n559_), .B1(new_n590_), .B2(new_n612_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT67), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT67), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n589_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT68), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n611_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n606_), .A2(new_n610_), .A3(KEYINPUT68), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(KEYINPUT12), .A3(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n625_), .B(new_n626_), .C1(new_n630_), .C2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n623_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT5), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT69), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT13), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n623_), .A2(new_n635_), .A3(new_n640_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n645_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT13), .B1(new_n642_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT70), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G232gat), .A2(G233gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT34), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT35), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n652_), .A2(KEYINPUT35), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT15), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n549_), .B(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n630_), .B2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n617_), .A2(new_n549_), .A3(new_n618_), .A4(new_n588_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT72), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n655_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G190gat), .B(G218gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(G134gat), .B(G162gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(KEYINPUT36), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n578_), .A2(new_n579_), .A3(new_n627_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT67), .B1(new_n617_), .B2(new_n618_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n588_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n550_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n590_), .A2(new_n662_), .A3(new_n549_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n661_), .A2(KEYINPUT72), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n655_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n672_), .A2(new_n675_), .A3(new_n676_), .A4(new_n657_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n664_), .A2(new_n668_), .A3(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n667_), .B(KEYINPUT36), .Z(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n664_), .B2(new_n677_), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n678_), .A2(new_n681_), .A3(KEYINPUT37), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT37), .B1(new_n678_), .B2(new_n681_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT76), .ZN(new_n687_));
  XNOR2_X1  g486(.A(G127gat), .B(G155gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(G183gat), .B(G211gat), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n689_), .B(new_n690_), .Z(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(KEYINPUT68), .A3(KEYINPUT17), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(KEYINPUT17), .B2(new_n691_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(G231gat), .A2(G233gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n611_), .B(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n521_), .A2(new_n524_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n693_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n697_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n692_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n685_), .A2(new_n702_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n558_), .A2(new_n650_), .A3(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n511_), .A3(new_n464_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT38), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n649_), .B(KEYINPUT70), .Z(new_n708_));
  NOR3_X1   g507(.A1(new_n708_), .A2(new_n557_), .A3(new_n702_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT98), .B1(new_n678_), .B2(new_n681_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n664_), .A2(new_n677_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n679_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT98), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n664_), .A2(new_n677_), .A3(new_n668_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n710_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n503_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n709_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G1gat), .B1(new_n719_), .B2(new_n483_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n705_), .A2(new_n706_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n707_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT99), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT99), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n707_), .A2(new_n724_), .A3(new_n720_), .A4(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1324gat));
  NAND3_X1  g525(.A1(new_n709_), .A2(new_n718_), .A3(new_n478_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G8gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT100), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(new_n730_), .A3(G8gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n729_), .A2(new_n731_), .A3(KEYINPUT39), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n727_), .B2(G8gat), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT39), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n321_), .A2(G8gat), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n733_), .A2(new_n734_), .B1(new_n704_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n732_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1325gat));
  OAI21_X1  g538(.A(G15gat), .B1(new_n719_), .B2(new_n502_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT41), .Z(new_n741_));
  XNOR2_X1  g540(.A(new_n500_), .B(KEYINPUT82), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n704_), .A2(new_n412_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1326gat));
  NAND3_X1  g543(.A1(new_n704_), .A2(new_n517_), .A3(new_n480_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G22gat), .B1(new_n719_), .B2(new_n405_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n746_), .A2(KEYINPUT103), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(KEYINPUT103), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n749_));
  AND3_X1   g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n745_), .B1(new_n750_), .B2(new_n751_), .ZN(G1327gat));
  NAND2_X1  g551(.A1(new_n717_), .A2(new_n702_), .ZN(new_n753_));
  NOR4_X1   g552(.A1(new_n503_), .A2(new_n708_), .A3(new_n557_), .A4(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G29gat), .B1(new_n754_), .B2(new_n464_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n480_), .A2(new_n321_), .A3(new_n483_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n489_), .A2(new_n305_), .A3(new_n318_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT33), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n760_), .A3(new_n492_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n494_), .B1(new_n294_), .B2(new_n300_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n495_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n762_), .B(new_n763_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n466_), .A2(new_n757_), .B1(new_n765_), .B2(new_n405_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n742_), .B1(new_n766_), .B2(new_n484_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n756_), .B(new_n685_), .C1(new_n767_), .C2(new_n465_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n503_), .B2(new_n684_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n650_), .A2(new_n556_), .A3(new_n702_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT44), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n774_), .B(new_n771_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n483_), .A2(new_n526_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n755_), .B1(new_n776_), .B2(new_n777_), .ZN(G1328gat));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n528_), .B1(new_n776_), .B2(new_n478_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n754_), .A2(new_n528_), .A3(new_n478_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n781_), .B(KEYINPUT45), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n773_), .A2(new_n775_), .A3(new_n321_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n785_), .B(KEYINPUT46), .C1(new_n786_), .C2(new_n528_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(G1329gat));
  INV_X1    g587(.A(G43gat), .ZN(new_n789_));
  NOR4_X1   g588(.A1(new_n773_), .A2(new_n775_), .A3(new_n789_), .A4(new_n440_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G43gat), .B1(new_n754_), .B2(new_n742_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT47), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n440_), .A2(new_n789_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n776_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(G1330gat));
  AOI21_X1  g596(.A(G50gat), .B1(new_n754_), .B2(new_n480_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n480_), .A2(G50gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n776_), .B2(new_n799_), .ZN(G1331gat));
  NOR2_X1   g599(.A1(new_n503_), .A2(new_n556_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n708_), .A2(KEYINPUT104), .A3(new_n703_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT104), .B1(new_n708_), .B2(new_n703_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n464_), .B1(new_n805_), .B2(KEYINPUT105), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT105), .ZN(new_n807_));
  NOR4_X1   g606(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .A4(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n602_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT106), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT106), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n602_), .C1(new_n806_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n701_), .A2(new_n557_), .ZN(new_n813_));
  NOR4_X1   g612(.A1(new_n503_), .A2(new_n650_), .A3(new_n717_), .A4(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n483_), .A2(new_n602_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n810_), .A2(new_n812_), .B1(new_n814_), .B2(new_n815_), .ZN(G1332gat));
  AOI21_X1  g615(.A(new_n600_), .B1(new_n814_), .B2(new_n478_), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT48), .Z(new_n818_));
  NAND3_X1  g617(.A1(new_n805_), .A2(new_n600_), .A3(new_n478_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1333gat));
  AOI21_X1  g619(.A(new_n592_), .B1(new_n814_), .B2(new_n742_), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n821_), .B(KEYINPUT49), .Z(new_n822_));
  NAND3_X1  g621(.A1(new_n805_), .A2(new_n592_), .A3(new_n742_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1334gat));
  AOI21_X1  g623(.A(new_n598_), .B1(new_n814_), .B2(new_n480_), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(KEYINPUT50), .Z(new_n826_));
  NAND3_X1  g625(.A1(new_n805_), .A2(new_n598_), .A3(new_n480_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(G1335gat));
  NOR2_X1   g627(.A1(new_n650_), .A2(new_n753_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n801_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT107), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT107), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n801_), .A2(new_n832_), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G85gat), .B1(new_n834_), .B2(new_n464_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n708_), .A2(new_n557_), .A3(new_n702_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n464_), .A2(G85gat), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT108), .Z(new_n839_));
  AOI21_X1  g638(.A(new_n835_), .B1(new_n837_), .B2(new_n839_), .ZN(G1336gat));
  INV_X1    g639(.A(G92gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n834_), .A2(new_n841_), .A3(new_n478_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n837_), .A2(new_n478_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT109), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1337gat));
  AOI21_X1  g645(.A(new_n562_), .B1(new_n837_), .B2(new_n742_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n500_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n834_), .B2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n849_), .B(new_n851_), .ZN(G1338gat));
  NAND3_X1  g651(.A1(new_n834_), .A2(new_n563_), .A3(new_n480_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n837_), .A2(new_n480_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(G106gat), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT52), .B(new_n563_), .C1(new_n837_), .C2(new_n480_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT53), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n860_), .B(new_n853_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1339gat));
  AND3_X1   g661(.A1(new_n548_), .A2(new_n552_), .A3(new_n506_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n645_), .B1(new_n863_), .B2(new_n553_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n625_), .B1(new_n630_), .B2(new_n634_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n559_), .B1(new_n865_), .B2(new_n621_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n635_), .A2(new_n867_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n632_), .A2(KEYINPUT12), .A3(new_n633_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n671_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n870_), .A2(KEYINPUT55), .A3(new_n625_), .A4(new_n626_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n866_), .A2(new_n868_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n641_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n872_), .A2(KEYINPUT56), .A3(new_n873_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n864_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n543_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n542_), .A2(new_n546_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n506_), .B1(new_n551_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n555_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n716_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n716_), .B(KEYINPUT57), .C1(new_n878_), .C2(new_n884_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n883_), .A2(new_n647_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n872_), .A2(KEYINPUT56), .A3(new_n873_), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT56), .B1(new_n872_), .B2(new_n873_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(KEYINPUT111), .A2(KEYINPUT58), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n889_), .B(new_n893_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n684_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n887_), .B(new_n888_), .C1(new_n897_), .C2(new_n898_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n897_), .A2(new_n898_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n702_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n813_), .B1(new_n648_), .B2(new_n646_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n684_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n902_), .A3(new_n684_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n901_), .A2(new_n907_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n406_), .A2(new_n440_), .A3(new_n483_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT59), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n909_), .B2(KEYINPUT115), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n913_), .B1(KEYINPUT115), .B2(new_n909_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n887_), .A2(new_n888_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n895_), .A2(new_n896_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n685_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n701_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n903_), .A2(new_n902_), .A3(new_n684_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n904_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n914_), .B1(new_n918_), .B2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT116), .B(G113gat), .Z(new_n922_));
  NAND4_X1  g721(.A1(new_n911_), .A2(new_n556_), .A3(new_n921_), .A4(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT113), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n910_), .A2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n909_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(new_n901_), .B2(new_n907_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT113), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n926_), .A2(new_n556_), .A3(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(G113gat), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT114), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(KEYINPUT114), .A3(new_n931_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n924_), .B1(new_n934_), .B2(new_n935_), .ZN(G1340gat));
  NAND2_X1  g735(.A1(new_n911_), .A2(new_n921_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT117), .B1(new_n937_), .B2(new_n650_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n911_), .A2(new_n939_), .A3(new_n708_), .A4(new_n921_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n938_), .A2(G120gat), .A3(new_n940_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n926_), .A2(new_n929_), .ZN(new_n942_));
  INV_X1    g741(.A(G120gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n650_), .B2(KEYINPUT60), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n942_), .B(new_n944_), .C1(KEYINPUT60), .C2(new_n943_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n941_), .A2(new_n945_), .ZN(G1341gat));
  NOR2_X1   g745(.A1(new_n702_), .A2(G127gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n926_), .A2(new_n929_), .A3(new_n947_), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n701_), .B(new_n921_), .C1(new_n928_), .C2(new_n912_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(G127gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(KEYINPUT118), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT118), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n948_), .A2(new_n950_), .A3(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n954_), .ZN(G1342gat));
  INV_X1    g754(.A(G134gat), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n942_), .A2(new_n956_), .A3(new_n717_), .ZN(new_n957_));
  OAI21_X1  g756(.A(G134gat), .B1(new_n937_), .B2(new_n684_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1343gat));
  NAND2_X1  g758(.A1(new_n917_), .A2(KEYINPUT112), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n897_), .A2(new_n898_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n915_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n920_), .B1(new_n962_), .B2(new_n702_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n502_), .A2(new_n480_), .ZN(new_n964_));
  NOR4_X1   g763(.A1(new_n963_), .A2(new_n478_), .A3(new_n483_), .A4(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(new_n556_), .ZN(new_n966_));
  XOR2_X1   g765(.A(KEYINPUT119), .B(G141gat), .Z(new_n967_));
  XNOR2_X1  g766(.A(new_n966_), .B(new_n967_), .ZN(G1344gat));
  NAND2_X1  g767(.A1(new_n965_), .A2(new_n708_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g769(.A1(new_n965_), .A2(new_n701_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(KEYINPUT61), .B(G155gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1346gat));
  AOI21_X1  g772(.A(G162gat), .B1(new_n965_), .B2(new_n717_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n685_), .A2(G162gat), .ZN(new_n975_));
  XOR2_X1   g774(.A(new_n975_), .B(KEYINPUT120), .Z(new_n976_));
  AOI21_X1  g775(.A(new_n974_), .B1(new_n965_), .B2(new_n976_), .ZN(G1347gat));
  NOR2_X1   g776(.A1(new_n918_), .A2(new_n920_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n478_), .A2(new_n483_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n502_), .A2(new_n979_), .ZN(new_n980_));
  INV_X1    g779(.A(new_n980_), .ZN(new_n981_));
  NOR3_X1   g780(.A1(new_n978_), .A2(new_n480_), .A3(new_n981_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(new_n556_), .ZN(new_n983_));
  OAI211_X1 g782(.A(KEYINPUT62), .B(G169gat), .C1(new_n983_), .C2(KEYINPUT22), .ZN(new_n984_));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n985_));
  INV_X1    g784(.A(new_n983_), .ZN(new_n986_));
  INV_X1    g785(.A(KEYINPUT22), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n985_), .B1(new_n986_), .B2(new_n987_), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n224_), .B1(new_n986_), .B2(new_n985_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n984_), .B1(new_n988_), .B2(new_n989_), .ZN(G1348gat));
  AOI21_X1  g789(.A(G176gat), .B1(new_n982_), .B2(new_n708_), .ZN(new_n991_));
  OAI21_X1  g790(.A(KEYINPUT121), .B1(new_n963_), .B2(new_n480_), .ZN(new_n992_));
  INV_X1    g791(.A(KEYINPUT121), .ZN(new_n993_));
  NAND3_X1  g792(.A1(new_n908_), .A2(new_n993_), .A3(new_n405_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n992_), .A2(new_n994_), .ZN(new_n995_));
  NOR3_X1   g794(.A1(new_n981_), .A2(new_n225_), .A3(new_n650_), .ZN(new_n996_));
  AOI21_X1  g795(.A(new_n991_), .B1(new_n995_), .B2(new_n996_), .ZN(G1349gat));
  NOR2_X1   g796(.A1(new_n978_), .A2(new_n480_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n217_), .A2(new_n221_), .ZN(new_n999_));
  NOR2_X1   g798(.A1(new_n981_), .A2(new_n702_), .ZN(new_n1000_));
  NAND3_X1  g799(.A1(new_n998_), .A2(new_n999_), .A3(new_n1000_), .ZN(new_n1001_));
  INV_X1    g800(.A(new_n1000_), .ZN(new_n1002_));
  AOI21_X1  g801(.A(new_n1002_), .B1(new_n992_), .B2(new_n994_), .ZN(new_n1003_));
  OAI21_X1  g802(.A(new_n1001_), .B1(new_n1003_), .B2(G183gat), .ZN(new_n1004_));
  NAND2_X1  g803(.A1(new_n1004_), .A2(KEYINPUT122), .ZN(new_n1005_));
  INV_X1    g804(.A(KEYINPUT122), .ZN(new_n1006_));
  OAI211_X1 g805(.A(new_n1001_), .B(new_n1006_), .C1(new_n1003_), .C2(G183gat), .ZN(new_n1007_));
  NAND2_X1  g806(.A1(new_n1005_), .A2(new_n1007_), .ZN(G1350gat));
  INV_X1    g807(.A(new_n982_), .ZN(new_n1009_));
  OAI21_X1  g808(.A(G190gat), .B1(new_n1009_), .B2(new_n684_), .ZN(new_n1010_));
  NAND3_X1  g809(.A1(new_n982_), .A2(new_n218_), .A3(new_n717_), .ZN(new_n1011_));
  NAND2_X1  g810(.A1(new_n1010_), .A2(new_n1011_), .ZN(G1351gat));
  INV_X1    g811(.A(KEYINPUT124), .ZN(new_n1013_));
  NOR2_X1   g812(.A1(new_n964_), .A2(new_n979_), .ZN(new_n1014_));
  INV_X1    g813(.A(new_n1014_), .ZN(new_n1015_));
  AOI21_X1  g814(.A(new_n1015_), .B1(new_n901_), .B2(new_n907_), .ZN(new_n1016_));
  AOI211_X1 g815(.A(new_n1013_), .B(G197gat), .C1(new_n1016_), .C2(new_n556_), .ZN(new_n1017_));
  NAND3_X1  g816(.A1(new_n908_), .A2(new_n556_), .A3(new_n1014_), .ZN(new_n1018_));
  AOI21_X1  g817(.A(KEYINPUT124), .B1(new_n1018_), .B2(new_n263_), .ZN(new_n1019_));
  NOR2_X1   g818(.A1(new_n1017_), .A2(new_n1019_), .ZN(new_n1020_));
  NAND4_X1  g819(.A1(new_n908_), .A2(G197gat), .A3(new_n556_), .A4(new_n1014_), .ZN(new_n1021_));
  NAND2_X1  g820(.A1(new_n1021_), .A2(KEYINPUT123), .ZN(new_n1022_));
  INV_X1    g821(.A(KEYINPUT123), .ZN(new_n1023_));
  NAND4_X1  g822(.A1(new_n1016_), .A2(new_n1023_), .A3(G197gat), .A4(new_n556_), .ZN(new_n1024_));
  AND2_X1   g823(.A1(new_n1022_), .A2(new_n1024_), .ZN(new_n1025_));
  OAI21_X1  g824(.A(KEYINPUT125), .B1(new_n1020_), .B2(new_n1025_), .ZN(new_n1026_));
  NAND2_X1  g825(.A1(new_n1022_), .A2(new_n1024_), .ZN(new_n1027_));
  INV_X1    g826(.A(KEYINPUT125), .ZN(new_n1028_));
  OAI211_X1 g827(.A(new_n1027_), .B(new_n1028_), .C1(new_n1019_), .C2(new_n1017_), .ZN(new_n1029_));
  NAND2_X1  g828(.A1(new_n1026_), .A2(new_n1029_), .ZN(G1352gat));
  NAND2_X1  g829(.A1(new_n1016_), .A2(new_n708_), .ZN(new_n1031_));
  XNOR2_X1  g830(.A(new_n1031_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g831(.A(new_n702_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1033_));
  NAND2_X1  g832(.A1(new_n1016_), .A2(new_n1033_), .ZN(new_n1034_));
  AND2_X1   g833(.A1(new_n1034_), .A2(KEYINPUT126), .ZN(new_n1035_));
  NOR2_X1   g834(.A1(new_n1034_), .A2(KEYINPUT126), .ZN(new_n1036_));
  NOR2_X1   g835(.A1(new_n1035_), .A2(new_n1036_), .ZN(new_n1037_));
  INV_X1    g836(.A(KEYINPUT63), .ZN(new_n1038_));
  NAND3_X1  g837(.A1(new_n1037_), .A2(new_n1038_), .A3(new_n255_), .ZN(new_n1039_));
  OAI22_X1  g838(.A1(new_n1035_), .A2(new_n1036_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1040_));
  NAND2_X1  g839(.A1(new_n1039_), .A2(new_n1040_), .ZN(G1354gat));
  NAND2_X1  g840(.A1(new_n1016_), .A2(new_n717_), .ZN(new_n1042_));
  XOR2_X1   g841(.A(KEYINPUT127), .B(G218gat), .Z(new_n1043_));
  NOR2_X1   g842(.A1(new_n684_), .A2(new_n1043_), .ZN(new_n1044_));
  AOI22_X1  g843(.A1(new_n1042_), .A2(new_n1043_), .B1(new_n1016_), .B2(new_n1044_), .ZN(G1355gat));
endmodule


