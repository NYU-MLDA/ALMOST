//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_, new_n977_,
    new_n978_, new_n979_, new_n981_, new_n982_, new_n983_, new_n985_,
    new_n986_, new_n987_, new_n989_, new_n990_, new_n991_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_, new_n999_;
  NOR2_X1   g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n204_), .B2(KEYINPUT9), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n203_), .A2(KEYINPUT65), .A3(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT65), .B1(new_n203_), .B2(new_n206_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n205_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT10), .B(G99gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT66), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n213_), .A2(new_n215_), .A3(G99gat), .A4(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n212_), .A2(KEYINPUT66), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n209_), .A2(new_n211_), .A3(new_n216_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n222_), .B(new_n223_), .C1(new_n224_), .C2(KEYINPUT67), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT67), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n224_), .A2(new_n222_), .A3(new_n223_), .A4(KEYINPUT67), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n220_), .A2(new_n227_), .A3(new_n216_), .A4(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n204_), .A2(new_n202_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n221_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT68), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G29gat), .B(G36gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G43gat), .B(G50gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(new_n221_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G232gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT35), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n238_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT15), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT15), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n238_), .A2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n252_), .A2(new_n234_), .B1(new_n245_), .B2(new_n244_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n241_), .A2(new_n247_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n247_), .B1(new_n241_), .B2(new_n253_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G190gat), .B(G218gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G134gat), .B(G162gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(KEYINPUT36), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n259_), .B(KEYINPUT36), .Z(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n264_), .A2(KEYINPUT37), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(KEYINPUT37), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G71gat), .B(G78gat), .Z(new_n268_));
  XNOR2_X1  g067(.A(G57gat), .B(G64gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(KEYINPUT11), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT69), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n268_), .B(new_n272_), .C1(KEYINPUT11), .C2(new_n269_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G15gat), .B(G22gat), .ZN(new_n279_));
  INV_X1    g078(.A(G1gat), .ZN(new_n280_));
  INV_X1    g079(.A(G8gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT14), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G1gat), .B(G8gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n284_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(G231gat), .B2(G233gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n278_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n287_), .B(new_n289_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n277_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n275_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G155gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT16), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G183gat), .B(G211gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT17), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n297_), .A2(new_n298_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT17), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n298_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n291_), .A2(new_n295_), .A3(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n291_), .A2(new_n295_), .B1(KEYINPUT17), .B2(new_n299_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT74), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n291_), .A2(new_n295_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n300_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n291_), .A2(new_n295_), .A3(new_n305_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n267_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n229_), .A2(new_n231_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT8), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n239_), .B1(new_n319_), .B2(new_n221_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n240_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n294_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n235_), .A2(new_n278_), .A3(new_n240_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(KEYINPUT70), .B(new_n294_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G230gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT64), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT12), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n322_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n278_), .A2(new_n332_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n234_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n331_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G120gat), .B(G148gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT5), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G176gat), .B(G204gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT71), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n329_), .A2(new_n336_), .A3(new_n342_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n347_));
  OR2_X1    g146(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n344_), .A2(KEYINPUT72), .A3(KEYINPUT13), .A4(new_n345_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n315_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT75), .ZN(new_n353_));
  OR2_X1    g152(.A1(G197gat), .A2(G204gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT21), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(KEYINPUT21), .A3(new_n355_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n359_), .A2(new_n360_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT78), .B(G176gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G169gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT23), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(G183gat), .A3(G190gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT89), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n372_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT89), .ZN(new_n377_));
  INV_X1    g176(.A(new_n374_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n368_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n367_), .A2(KEYINPUT24), .ZN(new_n382_));
  OR2_X1    g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT25), .B(G183gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT26), .B(G190gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n369_), .B2(KEYINPUT23), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n376_), .B2(new_n389_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n363_), .B1(new_n380_), .B2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n361_), .A2(new_n362_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n364_), .A2(new_n365_), .B1(G169gat), .B2(G176gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n391_), .B2(new_n374_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n387_), .A2(KEYINPUT77), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n385_), .A2(new_n386_), .A3(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n397_), .A2(new_n376_), .A3(new_n384_), .A4(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(new_n396_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n393_), .A2(new_n401_), .A3(KEYINPUT20), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n379_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n377_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n395_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n394_), .B(new_n408_), .C1(new_n391_), .C2(new_n388_), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n400_), .A2(new_n396_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n363_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n404_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n405_), .B1(new_n415_), .B2(KEYINPUT95), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(KEYINPUT95), .B2(new_n415_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT18), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n404_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n409_), .A2(new_n413_), .A3(KEYINPUT20), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n421_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT90), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n402_), .A2(new_n426_), .A3(new_n404_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n424_), .B(new_n425_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT27), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n424_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n421_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n429_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n422_), .A2(new_n432_), .B1(new_n435_), .B2(new_n431_), .ZN(new_n436_));
  INV_X1    g235(.A(G141gat), .ZN(new_n437_));
  INV_X1    g236(.A(G148gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT3), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(G141gat), .B2(G148gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G141gat), .A2(G148gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT2), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT82), .ZN(new_n446_));
  INV_X1    g245(.A(new_n443_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT2), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT82), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n442_), .A2(new_n446_), .A3(new_n448_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n453_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(KEYINPUT1), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT1), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(G155gat), .A3(G162gat), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n459_), .B(new_n461_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G141gat), .A2(G148gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n447_), .A2(new_n463_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n452_), .A2(new_n458_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT85), .B(KEYINPUT29), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT86), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n468_));
  INV_X1    g267(.A(new_n466_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n446_), .A2(new_n451_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n439_), .A2(new_n441_), .B1(new_n447_), .B2(KEYINPUT2), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n457_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n462_), .A2(new_n464_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n468_), .B(new_n469_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n467_), .A2(new_n474_), .A3(new_n363_), .ZN(new_n475_));
  INV_X1    g274(.A(G228gat), .ZN(new_n476_));
  INV_X1    g275(.A(G233gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT29), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n465_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n480_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n483_), .B(KEYINPUT84), .C1(new_n465_), .C2(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G78gat), .B(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n479_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n479_), .B2(new_n487_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G22gat), .B(G50gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT28), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n465_), .A2(new_n494_), .A3(new_n481_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n465_), .B2(new_n481_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n493_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n465_), .A2(new_n481_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT28), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n465_), .A2(new_n494_), .A3(new_n481_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n492_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n501_), .A3(KEYINPUT83), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT83), .B1(new_n497_), .B2(new_n501_), .ZN(new_n504_));
  OAI22_X1  g303(.A1(new_n490_), .A2(new_n491_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT87), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n479_), .A2(new_n487_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n488_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n478_), .A2(new_n475_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n489_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT87), .ZN(new_n512_));
  INV_X1    g311(.A(new_n504_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n502_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n511_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n491_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n497_), .A2(new_n501_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n509_), .B2(new_n489_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT88), .B1(new_n509_), .B2(new_n489_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n506_), .A2(new_n515_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G71gat), .B(G99gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G43gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n412_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G134gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G127gat), .ZN(new_n527_));
  INV_X1    g326(.A(G127gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G134gat), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT80), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n529_), .A3(KEYINPUT80), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G113gat), .B(G120gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n532_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n530_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n525_), .B(new_n538_), .Z(new_n539_));
  NAND2_X1  g338(.A1(G227gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(G15gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT30), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT31), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n539_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G225gat), .A2(G233gat), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n534_), .B(new_n537_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n538_), .A2(new_n465_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(KEYINPUT4), .ZN(new_n550_));
  OR3_X1    g349(.A1(new_n538_), .A2(new_n465_), .A3(KEYINPUT4), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n547_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G1gat), .B(G29gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(G85gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT0), .B(G57gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  INV_X1    g355(.A(new_n547_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n558_));
  OR3_X1    g357(.A1(new_n552_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n556_), .B1(new_n552_), .B2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n545_), .A2(new_n546_), .A3(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n436_), .A2(new_n522_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT97), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n417_), .A2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n433_), .A2(new_n566_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n561_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n550_), .A2(new_n551_), .A3(new_n547_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n556_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n548_), .A2(new_n549_), .A3(new_n557_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT93), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n550_), .A2(new_n551_), .A3(new_n547_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n574_), .A2(new_n577_), .B1(new_n560_), .B2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT33), .B(new_n556_), .C1(new_n552_), .C2(new_n558_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(KEYINPUT92), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(KEYINPUT92), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT91), .B1(new_n434_), .B2(new_n429_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n434_), .A2(KEYINPUT91), .A3(new_n429_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n569_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n517_), .A2(new_n521_), .A3(new_n519_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n505_), .A2(KEYINPUT87), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n512_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT96), .B1(new_n587_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n402_), .A2(new_n404_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT90), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n402_), .A2(new_n426_), .A3(new_n404_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n425_), .B1(new_n597_), .B2(new_n424_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n593_), .B1(new_n598_), .B2(new_n430_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n580_), .B(KEYINPUT92), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n599_), .A2(new_n586_), .A3(new_n600_), .A4(new_n579_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n567_), .A2(new_n568_), .A3(new_n561_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n591_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n561_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n436_), .A2(new_n591_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n592_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n545_), .A2(new_n546_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n565_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT76), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n249_), .A2(new_n287_), .A3(new_n251_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n238_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n287_), .A2(new_n248_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n614_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G169gat), .B(G197gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(new_n622_), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n616_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n616_), .B2(new_n620_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n612_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(KEYINPUT76), .A3(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n353_), .A2(new_n611_), .A3(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n280_), .A3(new_n561_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n264_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n611_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n349_), .A2(new_n350_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(new_n631_), .A3(new_n314_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n280_), .B1(new_n640_), .B2(new_n561_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n635_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n634_), .B2(new_n633_), .ZN(G1324gat));
  XNOR2_X1  g442(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n432_), .A2(new_n422_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n435_), .A2(new_n431_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n640_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT39), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n632_), .A2(new_n281_), .A3(new_n647_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n644_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n649_), .A2(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n648_), .B2(G8gat), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n651_), .B(new_n644_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n652_), .A2(new_n657_), .ZN(G1325gat));
  NAND3_X1  g457(.A1(new_n632_), .A2(new_n541_), .A3(new_n609_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n640_), .A2(new_n609_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(new_n660_), .B2(G15gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n522_), .B(KEYINPUT100), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n640_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n632_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n351_), .A2(new_n630_), .A3(new_n314_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT102), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  INV_X1    g477(.A(new_n267_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n607_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT96), .B(new_n591_), .C1(new_n602_), .C2(new_n601_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n610_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n565_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n678_), .B1(new_n684_), .B2(KEYINPUT103), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n686_), .B(KEYINPUT43), .C1(new_n611_), .C2(new_n679_), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n675_), .B(new_n677_), .C1(new_n685_), .C2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n561_), .A2(G29gat), .ZN(new_n689_));
  INV_X1    g488(.A(new_n677_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n682_), .A2(new_n683_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n267_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT43), .B1(new_n692_), .B2(new_n686_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n684_), .A2(KEYINPUT103), .A3(new_n678_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n675_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n677_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT104), .B1(new_n698_), .B2(KEYINPUT44), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n688_), .B(new_n689_), .C1(new_n697_), .C2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n611_), .A2(new_n631_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n308_), .A2(new_n313_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n264_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n638_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n701_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n561_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n674_), .B1(new_n700_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n707_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n697_), .A2(new_n699_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n698_), .A2(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT105), .B(new_n709_), .C1(new_n712_), .C2(new_n689_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n708_), .A2(new_n713_), .ZN(G1328gat));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  INV_X1    g514(.A(G36gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n688_), .A2(new_n436_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n710_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n647_), .A2(KEYINPUT106), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n647_), .A2(KEYINPUT106), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n720_), .B1(new_n706_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n701_), .A2(new_n705_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n725_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n727_), .A2(KEYINPUT107), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n719_), .B1(new_n726_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n706_), .A2(new_n720_), .A3(new_n725_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT107), .B1(new_n727_), .B2(new_n728_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(KEYINPUT45), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n715_), .B1(new_n718_), .B2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n730_), .A2(new_n733_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n711_), .A2(new_n647_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n699_), .B2(new_n697_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n736_), .B(KEYINPUT46), .C1(new_n738_), .C2(new_n716_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n735_), .A2(new_n739_), .ZN(G1329gat));
  NAND2_X1  g539(.A1(new_n609_), .A2(G43gat), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n688_), .B(new_n741_), .C1(new_n697_), .C2(new_n699_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G43gat), .B1(new_n706_), .B2(new_n609_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT47), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745_));
  INV_X1    g544(.A(new_n743_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n745_), .B(new_n746_), .C1(new_n712_), .C2(new_n741_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(G1330gat));
  INV_X1    g547(.A(G50gat), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n688_), .A2(new_n522_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n710_), .B2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n667_), .A2(G50gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT108), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n706_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT109), .B1(new_n751_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n711_), .A2(new_n591_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n699_), .B2(new_n697_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n757_), .B(new_n754_), .C1(new_n759_), .C2(new_n749_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n756_), .A2(new_n760_), .ZN(G1331gat));
  NOR2_X1   g560(.A1(new_n611_), .A2(new_n630_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n762_), .A2(new_n638_), .A3(new_n315_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G57gat), .B1(new_n763_), .B2(new_n561_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT110), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n351_), .A2(new_n630_), .A3(new_n314_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n637_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT111), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n637_), .A2(new_n769_), .A3(new_n766_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n561_), .A2(G57gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n765_), .B1(new_n771_), .B2(new_n772_), .ZN(G1332gat));
  INV_X1    g572(.A(G64gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n763_), .A2(new_n774_), .A3(new_n723_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n768_), .A2(new_n723_), .A3(new_n770_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(G64gat), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G64gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT113), .B(new_n775_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1333gat));
  INV_X1    g583(.A(G71gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n763_), .A2(new_n785_), .A3(new_n609_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n771_), .A2(new_n609_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G71gat), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(KEYINPUT49), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(KEYINPUT49), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1334gat));
  INV_X1    g590(.A(G78gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n763_), .A2(new_n792_), .A3(new_n668_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n771_), .A2(new_n668_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G78gat), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(KEYINPUT50), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(KEYINPUT50), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(G1335gat));
  NOR3_X1   g597(.A1(new_n351_), .A2(new_n630_), .A3(new_n702_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806_), .B2(new_n606_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n351_), .A2(new_n704_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n762_), .A2(new_n808_), .ZN(new_n809_));
  OR3_X1    g608(.A1(new_n809_), .A2(G85gat), .A3(new_n606_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(G1336gat));
  OAI21_X1  g610(.A(G92gat), .B1(new_n806_), .B2(new_n724_), .ZN(new_n812_));
  OR3_X1    g611(.A1(new_n809_), .A2(G92gat), .A3(new_n436_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1337gat));
  NOR3_X1   g613(.A1(new_n809_), .A2(new_n610_), .A3(new_n210_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n610_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n222_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT51), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n816_), .C1(new_n817_), .C2(new_n222_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1338gat));
  NAND4_X1  g621(.A1(new_n762_), .A2(new_n223_), .A3(new_n591_), .A4(new_n808_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n801_), .A2(new_n591_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(G106gat), .ZN(new_n826_));
  AOI211_X1 g625(.A(KEYINPUT52), .B(new_n223_), .C1(new_n801_), .C2(new_n591_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n278_), .B1(new_n235_), .B2(new_n240_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n335_), .B1(new_n833_), .B2(KEYINPUT12), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n324_), .A2(new_n330_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT55), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n331_), .A2(new_n333_), .A3(new_n837_), .A4(new_n335_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n333_), .A2(new_n335_), .A3(new_n324_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n836_), .A2(new_n838_), .B1(new_n839_), .B2(new_n328_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n341_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n832_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n832_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n839_), .A2(new_n328_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n322_), .A2(new_n332_), .B1(new_n234_), .B2(new_n334_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n837_), .B1(new_n848_), .B2(new_n331_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n834_), .A2(KEYINPUT55), .A3(new_n835_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(KEYINPUT116), .A3(new_n844_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n842_), .A2(new_n846_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n329_), .A2(new_n336_), .A3(new_n841_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n854_), .A2(new_n630_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n613_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n623_), .B1(new_n618_), .B2(new_n615_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n625_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n346_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(KEYINPUT57), .A3(new_n264_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n860_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n636_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n851_), .A2(new_n844_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n842_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT117), .B1(new_n854_), .B2(new_n859_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n854_), .A2(KEYINPUT117), .A3(new_n859_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n867_), .B1(new_n869_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n842_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n875_), .A2(KEYINPUT58), .A3(new_n872_), .A4(new_n871_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n876_), .A3(new_n267_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n863_), .A2(new_n866_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n314_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n314_), .B2(new_n630_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n631_), .A2(new_n702_), .A3(KEYINPUT115), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n266_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n264_), .A2(KEYINPUT37), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n351_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n882_), .B(new_n881_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT54), .B1(new_n889_), .B2(new_n638_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n831_), .B1(new_n879_), .B2(new_n892_), .ZN(new_n893_));
  AOI211_X1 g692(.A(KEYINPUT118), .B(new_n891_), .C1(new_n878_), .C2(new_n314_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n647_), .A2(new_n591_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n610_), .A2(new_n606_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n830_), .B1(new_n895_), .B2(new_n899_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n865_), .A2(new_n864_), .A3(new_n636_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n866_), .A2(new_n877_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n866_), .A2(new_n877_), .A3(KEYINPUT119), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n702_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n830_), .B(new_n899_), .C1(new_n906_), .C2(new_n891_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT120), .B1(new_n900_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n893_), .A2(new_n894_), .A3(new_n898_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n910_), .B(new_n907_), .C1(new_n911_), .C2(new_n830_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n630_), .A2(G113gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT121), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n909_), .A2(new_n912_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(G113gat), .ZN(new_n916_));
  INV_X1    g715(.A(new_n911_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n631_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n915_), .A2(new_n918_), .ZN(G1340gat));
  XOR2_X1   g718(.A(KEYINPUT122), .B(G120gat), .Z(new_n920_));
  NOR2_X1   g719(.A1(new_n351_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n911_), .B1(KEYINPUT60), .B2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n638_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n907_), .B1(new_n911_), .B2(new_n830_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n920_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(KEYINPUT60), .B2(new_n922_), .ZN(G1341gat));
  NOR2_X1   g725(.A1(new_n314_), .A2(new_n528_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n909_), .A2(new_n912_), .A3(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n893_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n894_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n929_), .A2(new_n930_), .A3(new_n702_), .A4(new_n899_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n931_), .A2(KEYINPUT123), .A3(new_n528_), .ZN(new_n932_));
  AOI21_X1  g731(.A(KEYINPUT123), .B1(new_n931_), .B2(new_n528_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n928_), .A2(new_n934_), .ZN(G1342gat));
  NOR2_X1   g734(.A1(new_n679_), .A2(new_n526_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n909_), .A2(new_n912_), .A3(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n526_), .B1(new_n917_), .B2(new_n264_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1343gat));
  NOR3_X1   g738(.A1(new_n723_), .A2(new_n522_), .A3(new_n606_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n895_), .A2(new_n610_), .A3(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n631_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n437_), .ZN(G1344gat));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n351_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(new_n438_), .ZN(G1345gat));
  OAI21_X1  g744(.A(KEYINPUT124), .B1(new_n941_), .B2(new_n314_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n893_), .A2(new_n894_), .A3(new_n609_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n947_), .A2(new_n948_), .A3(new_n702_), .A4(new_n940_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(KEYINPUT61), .B(G155gat), .ZN(new_n950_));
  AND3_X1   g749(.A1(new_n946_), .A2(new_n949_), .A3(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n946_), .B2(new_n949_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1346gat));
  OAI21_X1  g752(.A(G162gat), .B1(new_n941_), .B2(new_n679_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n264_), .A2(G162gat), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n941_), .B2(new_n955_), .ZN(G1347gat));
  NOR2_X1   g755(.A1(new_n906_), .A2(new_n891_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n723_), .A2(new_n562_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n959_), .A2(new_n630_), .A3(new_n667_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G169gat), .B1(new_n957_), .B2(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n957_), .A2(new_n960_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(new_n365_), .ZN(new_n965_));
  OAI211_X1 g764(.A(KEYINPUT62), .B(G169gat), .C1(new_n957_), .C2(new_n960_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n963_), .A2(new_n965_), .A3(new_n966_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n963_), .A2(new_n965_), .A3(KEYINPUT125), .A4(new_n966_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1348gat));
  NOR3_X1   g770(.A1(new_n957_), .A2(new_n668_), .A3(new_n958_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(new_n638_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n893_), .A2(new_n894_), .A3(new_n591_), .ZN(new_n974_));
  AND3_X1   g773(.A1(new_n959_), .A2(G176gat), .A3(new_n638_), .ZN(new_n975_));
  AOI22_X1  g774(.A1(new_n973_), .A2(new_n364_), .B1(new_n974_), .B2(new_n975_), .ZN(G1349gat));
  NAND3_X1  g775(.A1(new_n974_), .A2(new_n702_), .A3(new_n959_), .ZN(new_n977_));
  INV_X1    g776(.A(G183gat), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n314_), .A2(new_n385_), .ZN(new_n979_));
  AOI22_X1  g778(.A1(new_n977_), .A2(new_n978_), .B1(new_n972_), .B2(new_n979_), .ZN(G1350gat));
  NAND3_X1  g779(.A1(new_n972_), .A2(new_n386_), .A3(new_n636_), .ZN(new_n981_));
  AND2_X1   g780(.A1(new_n972_), .A2(new_n267_), .ZN(new_n982_));
  INV_X1    g781(.A(G190gat), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n981_), .B1(new_n982_), .B2(new_n983_), .ZN(G1351gat));
  NOR3_X1   g783(.A1(new_n724_), .A2(new_n522_), .A3(new_n561_), .ZN(new_n985_));
  AND2_X1   g784(.A1(new_n947_), .A2(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(new_n630_), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n987_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g787(.A1(new_n947_), .A2(new_n985_), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n989_), .A2(new_n351_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(KEYINPUT126), .B(G204gat), .ZN(new_n991_));
  XNOR2_X1  g790(.A(new_n990_), .B(new_n991_), .ZN(G1353gat));
  AOI21_X1  g791(.A(new_n314_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n986_), .A2(new_n993_), .ZN(new_n994_));
  OR2_X1    g793(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n994_), .B(new_n995_), .ZN(G1354gat));
  XOR2_X1   g795(.A(KEYINPUT127), .B(G218gat), .Z(new_n997_));
  NOR3_X1   g796(.A1(new_n989_), .A2(new_n679_), .A3(new_n997_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n986_), .A2(new_n636_), .ZN(new_n999_));
  AOI21_X1  g798(.A(new_n998_), .B1(new_n999_), .B2(new_n997_), .ZN(G1355gat));
endmodule


