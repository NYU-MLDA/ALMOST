//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G85gat), .B(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT10), .B(G99gat), .Z(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n211_), .A2(KEYINPUT9), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(new_n210_), .B2(KEYINPUT65), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT7), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n217_), .B(new_n211_), .C1(new_n205_), .C2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n211_), .B1(new_n205_), .B2(new_n222_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n217_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n215_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n235_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n209_), .A2(new_n214_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(new_n223_), .A3(new_n234_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n202_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n234_), .B1(new_n237_), .B2(new_n223_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT12), .B1(new_n242_), .B2(KEYINPUT67), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT67), .B1(new_n227_), .B2(new_n235_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n243_), .A2(new_n246_), .A3(new_n202_), .A4(new_n238_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n239_), .A2(new_n240_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G120gat), .B(G148gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT5), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G176gat), .B(G204gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n250_), .B(new_n251_), .Z(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n241_), .A2(new_n247_), .A3(new_n248_), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n239_), .B(KEYINPUT66), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n257_), .A2(KEYINPUT68), .A3(new_n247_), .A4(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n247_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n252_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT13), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT13), .B1(new_n259_), .B2(new_n261_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G229gat), .A2(G233gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT74), .B(G8gat), .Z(new_n269_));
  INV_X1    g068(.A(G1gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT14), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G15gat), .B(G22gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G1gat), .B(G8gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n273_), .B(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G29gat), .B(G36gat), .Z(new_n277_));
  XOR2_X1   g076(.A(G43gat), .B(G50gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n276_), .A2(new_n279_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n268_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n279_), .B(KEYINPUT15), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n273_), .B(new_n274_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(new_n267_), .A3(new_n280_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G141gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G169gat), .B(G197gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  AND3_X1   g090(.A1(new_n288_), .A2(KEYINPUT77), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n288_), .B2(KEYINPUT77), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n266_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT85), .ZN(new_n297_));
  INV_X1    g096(.A(G204gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G197gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G197gat), .A2(G204gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT21), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n303_), .B1(new_n301_), .B2(G197gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n309_), .B2(KEYINPUT21), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n298_), .A2(G197gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(G197gat), .B1(new_n299_), .B2(new_n300_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(KEYINPUT86), .ZN(new_n313_));
  INV_X1    g112(.A(G197gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(KEYINPUT86), .B(new_n314_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT21), .B1(new_n313_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n310_), .B1(new_n319_), .B2(KEYINPUT87), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT86), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n321_), .A2(new_n322_), .B1(G197gat), .B2(new_n298_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n306_), .B1(new_n323_), .B2(new_n317_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n308_), .B1(new_n320_), .B2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(KEYINPUT78), .B(G190gat), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT26), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(KEYINPUT26), .B2(G190gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT25), .B(G183gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT23), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G169gat), .ZN(new_n339_));
  INV_X1    g138(.A(G176gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n341_), .A2(new_n336_), .A3(new_n335_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n332_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n334_), .B1(G183gat), .B2(new_n328_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT22), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n339_), .B1(new_n347_), .B2(new_n340_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n335_), .B2(new_n347_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n296_), .B1(new_n327_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT91), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n338_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n331_), .B(KEYINPUT90), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G190gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n342_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT22), .B(G169gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n340_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT92), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n361_), .A2(new_n362_), .B1(new_n334_), .B2(new_n364_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n355_), .A2(new_n358_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n353_), .B1(new_n327_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT19), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n308_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n307_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n319_), .A2(KEYINPUT87), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n371_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n344_), .A2(new_n350_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(KEYINPUT93), .A3(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n352_), .A2(new_n367_), .A3(new_n370_), .A4(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT20), .B1(new_n376_), .B2(new_n377_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n327_), .A2(new_n366_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n369_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G8gat), .B(G36gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n379_), .A2(new_n382_), .A3(new_n388_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(KEYINPUT95), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT27), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT95), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n383_), .A2(new_n394_), .A3(new_n389_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G228gat), .ZN(new_n397_));
  INV_X1    g196(.A(G233gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G141gat), .A2(G148gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G155gat), .A2(G162gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(KEYINPUT1), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT1), .ZN(new_n410_));
  INV_X1    g209(.A(new_n407_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n409_), .A2(KEYINPUT81), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n413_), .B(new_n407_), .C1(new_n408_), .C2(KEYINPUT1), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n406_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n411_), .A2(new_n408_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT3), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n404_), .A2(KEYINPUT82), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n420_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n402_), .B(KEYINPUT2), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n417_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n401_), .B1(new_n415_), .B2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n402_), .B(KEYINPUT2), .Z(new_n427_));
  OAI21_X1  g226(.A(new_n416_), .B1(new_n427_), .B2(new_n422_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n409_), .A2(KEYINPUT81), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n411_), .A2(new_n410_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n429_), .A2(new_n414_), .A3(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT83), .B(new_n428_), .C1(new_n431_), .C2(new_n406_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n426_), .A2(new_n432_), .A3(KEYINPUT29), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n376_), .A2(new_n400_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT88), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n412_), .A2(new_n414_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n424_), .A2(new_n421_), .A3(new_n419_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n436_), .A2(new_n405_), .B1(new_n437_), .B2(new_n416_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n435_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT88), .B(KEYINPUT29), .C1(new_n415_), .C2(new_n425_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(KEYINPUT89), .B(new_n399_), .C1(new_n442_), .C2(new_n327_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n376_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT89), .B1(new_n445_), .B2(new_n399_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n434_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G78gat), .B(G106gat), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n426_), .A2(new_n432_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n439_), .ZN(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n439_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G22gat), .B(G50gat), .Z(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n457_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n459_), .A3(new_n455_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n399_), .B1(new_n442_), .B2(new_n327_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n443_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n448_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n434_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n449_), .A2(new_n462_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n466_), .B2(new_n434_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n434_), .ZN(new_n471_));
  AOI211_X1 g270(.A(new_n448_), .B(new_n471_), .C1(new_n465_), .C2(new_n443_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n461_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n380_), .A2(new_n381_), .A3(new_n369_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n352_), .A2(new_n367_), .A3(new_n378_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n369_), .B2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT27), .B(new_n391_), .C1(new_n476_), .C2(new_n388_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n396_), .A2(new_n469_), .A3(new_n473_), .A4(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT100), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n473_), .A2(new_n469_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT100), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n396_), .A4(new_n477_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT80), .B(G15gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n377_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G127gat), .B(G134gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G113gat), .B(G120gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n489_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n487_), .B(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G71gat), .B(G99gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(G43gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT30), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT31), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n493_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G225gat), .A2(G233gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n500_), .B(KEYINPUT98), .Z(new_n501_));
  NAND3_X1  g300(.A1(new_n426_), .A2(new_n432_), .A3(new_n492_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n492_), .A2(KEYINPUT96), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n490_), .A2(new_n491_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n438_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n501_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n502_), .A2(KEYINPUT4), .A3(new_n507_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT97), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n502_), .A2(new_n511_), .A3(new_n507_), .A4(KEYINPUT4), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n502_), .A2(KEYINPUT4), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n508_), .B1(new_n515_), .B2(new_n501_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G29gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G85gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT0), .B(G57gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n501_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n513_), .B1(KEYINPUT97), .B2(new_n509_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(new_n512_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n525_), .B2(new_n508_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n499_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n483_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n473_), .A2(new_n469_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n527_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n530_), .A2(new_n396_), .A3(new_n531_), .A4(new_n477_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n523_), .A3(new_n512_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n502_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n534_), .A2(new_n521_), .A3(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT33), .B1(new_n516_), .B2(new_n521_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT33), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n538_), .B(new_n520_), .C1(new_n525_), .C2(new_n508_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n392_), .A2(new_n395_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n388_), .A2(KEYINPUT32), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT99), .B1(new_n476_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT99), .ZN(new_n545_));
  INV_X1    g344(.A(new_n543_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n475_), .A2(new_n369_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n545_), .B(new_n546_), .C1(new_n547_), .C2(new_n474_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n379_), .A2(new_n382_), .A3(new_n543_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n527_), .A2(new_n544_), .A3(new_n548_), .A4(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n530_), .B1(new_n542_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n499_), .B1(new_n533_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n295_), .B1(new_n529_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT37), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(KEYINPUT37), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT70), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n562_), .B2(KEYINPUT72), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n284_), .A2(new_n227_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n237_), .A2(new_n223_), .A3(new_n279_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n562_), .A2(KEYINPUT72), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n569_), .A2(new_n563_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G190gat), .B(G218gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT71), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT36), .Z(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n570_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n574_), .A2(KEYINPUT36), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n555_), .B(new_n556_), .C1(new_n577_), .C2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n582_), .A2(new_n554_), .A3(KEYINPUT37), .A4(new_n576_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n234_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n285_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n588_), .A2(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n585_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT76), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n553_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n270_), .A3(new_n527_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n582_), .A2(new_n576_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(new_n598_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n553_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n531_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n604_), .A2(new_n605_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(new_n611_), .A3(new_n612_), .ZN(G1324gat));
  NAND2_X1  g412(.A1(new_n396_), .A2(new_n477_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n610_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT101), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n618_), .B(G8gat), .C1(new_n610_), .C2(new_n615_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(KEYINPUT39), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(KEYINPUT101), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n603_), .A2(new_n269_), .A3(new_n614_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT40), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n620_), .A2(KEYINPUT40), .A3(new_n622_), .A4(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(G1325gat));
  OAI21_X1  g427(.A(G15gat), .B1(new_n610_), .B2(new_n499_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT41), .Z(new_n630_));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n603_), .A2(new_n631_), .A3(new_n498_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(G1326gat));
  OAI21_X1  g432(.A(G22gat), .B1(new_n610_), .B2(new_n480_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n603_), .A2(new_n636_), .A3(new_n530_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1327gat));
  NOR2_X1   g437(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n584_), .B(KEYINPUT102), .Z(new_n640_));
  NAND2_X1  g439(.A1(new_n542_), .A2(new_n550_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n480_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n498_), .B1(new_n642_), .B2(new_n532_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n528_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n640_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n529_), .A2(new_n552_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n584_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n646_), .A2(KEYINPUT43), .B1(new_n647_), .B2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n295_), .A2(new_n599_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n639_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n639_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n648_), .B1(new_n647_), .B2(new_n640_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n649_), .B1(new_n529_), .B2(new_n552_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n652_), .B(new_n655_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(new_n527_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G29gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n295_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n607_), .A2(new_n599_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n661_), .B(new_n662_), .C1(new_n643_), .C2(new_n645_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n531_), .A2(G29gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n654_), .A2(new_n614_), .A3(new_n658_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n615_), .A2(G36gat), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT104), .B1(new_n663_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n553_), .A2(new_n671_), .A3(new_n662_), .A4(new_n668_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n670_), .A2(new_n672_), .A3(KEYINPUT45), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT45), .B1(new_n670_), .B2(new_n672_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n667_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n667_), .A2(KEYINPUT46), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1329gat));
  NOR3_X1   g479(.A1(new_n663_), .A2(G43gat), .A3(new_n499_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n654_), .A2(new_n498_), .A3(new_n658_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(G43gat), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n684_), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n681_), .B(new_n686_), .C1(new_n682_), .C2(G43gat), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1330gat));
  NAND3_X1  g487(.A1(new_n654_), .A2(new_n530_), .A3(new_n658_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G50gat), .ZN(new_n690_));
  OR3_X1    g489(.A1(new_n663_), .A2(G50gat), .A3(new_n480_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT106), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n690_), .A2(new_n694_), .A3(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1331gat));
  NOR2_X1   g495(.A1(new_n266_), .A2(new_n294_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n647_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n609_), .ZN(new_n699_));
  INV_X1    g498(.A(G57gat), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n531_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n602_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n531_), .B1(new_n702_), .B2(KEYINPUT107), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(KEYINPUT107), .B2(new_n702_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n701_), .B1(new_n704_), .B2(new_n700_), .ZN(G1332gat));
  NAND3_X1  g504(.A1(new_n698_), .A2(new_n614_), .A3(new_n609_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(G64gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n706_), .B2(G64gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n615_), .A2(G64gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT108), .Z(new_n712_));
  OAI22_X1  g511(.A1(new_n709_), .A2(new_n710_), .B1(new_n702_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT109), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715_));
  OAI221_X1 g514(.A(new_n715_), .B1(new_n702_), .B2(new_n712_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n699_), .B2(new_n499_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT49), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n499_), .A2(G71gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n702_), .B2(new_n720_), .ZN(G1334gat));
  OAI21_X1  g520(.A(G78gat), .B1(new_n699_), .B2(new_n480_), .ZN(new_n722_));
  XOR2_X1   g521(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n480_), .A2(G78gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n702_), .B2(new_n725_), .ZN(G1335gat));
  NAND2_X1  g525(.A1(new_n698_), .A2(new_n662_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G85gat), .B1(new_n728_), .B2(new_n527_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n646_), .A2(KEYINPUT43), .ZN(new_n730_));
  INV_X1    g529(.A(new_n657_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n697_), .A2(new_n598_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n527_), .A2(G85gat), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT112), .Z(new_n738_));
  AOI21_X1  g537(.A(new_n729_), .B1(new_n736_), .B2(new_n738_), .ZN(G1336gat));
  AOI21_X1  g538(.A(G92gat), .B1(new_n728_), .B2(new_n614_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n614_), .A2(new_n206_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n736_), .B2(new_n741_), .ZN(G1337gat));
  INV_X1    g541(.A(G99gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n736_), .B2(new_n498_), .ZN(new_n744_));
  AND4_X1   g543(.A1(new_n212_), .A2(new_n698_), .A3(new_n498_), .A4(new_n662_), .ZN(new_n745_));
  OR3_X1    g544(.A1(new_n744_), .A2(KEYINPUT51), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT51), .B1(new_n744_), .B2(new_n745_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1338gat));
  NAND3_X1  g547(.A1(new_n728_), .A2(new_n213_), .A3(new_n530_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n735_), .B(new_n530_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G106gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G106gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n749_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  NAND3_X1  g557(.A1(new_n483_), .A2(new_n527_), .A3(new_n498_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT116), .Z(new_n760_));
  NOR3_X1   g559(.A1(new_n584_), .A2(new_n294_), .A3(new_n598_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n266_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(new_n266_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  INV_X1    g565(.A(new_n291_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n281_), .A2(new_n282_), .A3(new_n268_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n267_), .B1(new_n286_), .B2(new_n280_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n283_), .A2(new_n287_), .A3(new_n291_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n294_), .A2(new_n259_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n202_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n246_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n238_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(KEYINPUT55), .ZN(new_n779_));
  INV_X1    g578(.A(new_n777_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n780_), .A2(KEYINPUT113), .A3(new_n202_), .A4(new_n246_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n247_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n779_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n778_), .A2(KEYINPUT55), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n783_), .A3(new_n781_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n253_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n774_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n788_), .A2(new_n789_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n773_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n766_), .B1(new_n792_), .B2(new_n608_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n773_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n788_), .A2(new_n789_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n774_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n788_), .A2(new_n789_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT57), .A3(new_n607_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(KEYINPUT58), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n788_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n772_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n788_), .B2(new_n803_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n802_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n788_), .A2(new_n803_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n802_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n804_), .A4(new_n806_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n811_), .A3(new_n584_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n793_), .A2(new_n800_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n765_), .B1(new_n813_), .B2(new_n598_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n760_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n294_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n294_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n815_), .A2(KEYINPUT59), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(KEYINPUT59), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n821_), .B2(new_n816_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n266_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n815_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n266_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n823_), .ZN(G1341gat));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n815_), .A2(new_n828_), .A3(new_n599_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n598_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n828_), .ZN(G1342gat));
  NAND2_X1  g630(.A1(new_n584_), .A2(G134gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n833_));
  AOI211_X1 g632(.A(KEYINPUT117), .B(G134gat), .C1(new_n815_), .C2(new_n608_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G134gat), .B1(new_n815_), .B2(new_n608_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n833_), .A2(new_n834_), .A3(new_n837_), .ZN(G1343gat));
  INV_X1    g637(.A(new_n814_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n614_), .A2(new_n480_), .A3(new_n531_), .A4(new_n498_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n818_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT118), .B(G141gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  INV_X1    g643(.A(new_n841_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n266_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g647(.A1(new_n841_), .A2(KEYINPUT119), .A3(new_n598_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT119), .B1(new_n841_), .B2(new_n598_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1346gat));
  AOI21_X1  g653(.A(G162gat), .B1(new_n845_), .B2(new_n608_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n640_), .A2(G162gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n845_), .B2(new_n856_), .ZN(G1347gat));
  NOR2_X1   g656(.A1(new_n644_), .A2(new_n530_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n814_), .A2(new_n615_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n294_), .A2(new_n359_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT121), .Z(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n814_), .A2(new_n818_), .A3(new_n615_), .A4(new_n859_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n339_), .B1(new_n864_), .B2(KEYINPUT120), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n814_), .A2(new_n615_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n294_), .A3(new_n858_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n865_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n865_), .B2(new_n869_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n863_), .B1(new_n871_), .B2(new_n872_), .ZN(G1348gat));
  INV_X1    g672(.A(new_n860_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n340_), .B1(new_n874_), .B2(new_n266_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT122), .B(new_n340_), .C1(new_n874_), .C2(new_n266_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n860_), .A2(G176gat), .A3(new_n846_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n880_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n877_), .A2(new_n878_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  NAND2_X1  g682(.A1(new_n860_), .A2(new_n599_), .ZN(new_n884_));
  MUX2_X1   g683(.A(new_n356_), .B(G183gat), .S(new_n884_), .Z(G1350gat));
  OAI21_X1  g684(.A(G190gat), .B1(new_n874_), .B2(new_n585_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n860_), .A2(new_n357_), .A3(new_n608_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1351gat));
  NAND3_X1  g687(.A1(new_n530_), .A2(new_n499_), .A3(new_n531_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT124), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n866_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n818_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n314_), .ZN(G1352gat));
  AND3_X1   g692(.A1(new_n839_), .A2(new_n614_), .A3(new_n890_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n846_), .A3(new_n301_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n298_), .B1(new_n891_), .B2(new_n266_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1353gat));
  INV_X1    g699(.A(KEYINPUT127), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n598_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT126), .Z(new_n903_));
  AND3_X1   g702(.A1(new_n894_), .A2(new_n901_), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n901_), .B1(new_n894_), .B2(new_n903_), .ZN(new_n905_));
  OAI22_X1  g704(.A1(new_n904_), .A2(new_n905_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n894_), .A2(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT127), .ZN(new_n908_));
  NOR2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n894_), .A2(new_n901_), .A3(new_n903_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n906_), .A2(new_n911_), .ZN(G1354gat));
  OR3_X1    g711(.A1(new_n891_), .A2(G218gat), .A3(new_n607_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G218gat), .B1(new_n891_), .B2(new_n585_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1355gat));
endmodule


