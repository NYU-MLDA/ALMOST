//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_;
  XOR2_X1   g000(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT78), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G134gat), .B(G162gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT79), .B(KEYINPUT36), .Z(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G85gat), .B(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT67), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT6), .ZN(new_n219_));
  INV_X1    g018(.A(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI22_X1  g021(.A1(new_n217_), .A2(new_n219_), .B1(KEYINPUT7), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n213_), .B1(new_n215_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT8), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(new_n213_), .C1(new_n215_), .C2(new_n223_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n229_), .A2(KEYINPUT64), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT64), .B1(new_n229_), .B2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n221_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n234_));
  INV_X1    g033(.A(G85gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n238_), .B2(KEYINPUT9), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n217_), .A2(new_n219_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT66), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n233_), .A2(new_n239_), .A3(new_n243_), .A4(new_n240_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n245_), .A2(KEYINPUT74), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(KEYINPUT74), .ZN(new_n247_));
  XOR2_X1   g046(.A(G43gat), .B(G50gat), .Z(new_n248_));
  OR3_X1    g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n228_), .A2(new_n242_), .A3(new_n244_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT34), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT35), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(KEYINPUT35), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT73), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n251_), .B(KEYINPUT15), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n228_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT76), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n255_), .B2(new_n260_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n252_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT75), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n271_), .A2(KEYINPUT76), .A3(new_n254_), .A4(new_n259_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n264_), .A2(new_n265_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(KEYINPUT77), .A3(new_n263_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT77), .B1(new_n274_), .B2(new_n263_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n211_), .B(new_n267_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n267_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n277_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n275_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n207_), .B(KEYINPUT36), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT37), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G57gat), .B(G64gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n286_));
  XOR2_X1   g085(.A(G71gat), .B(G78gat), .Z(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n265_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT71), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n296_), .A3(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G230gat), .A2(G233gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n265_), .A2(new_n291_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n265_), .A2(KEYINPUT12), .A3(new_n291_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n265_), .A2(KEYINPUT69), .A3(KEYINPUT12), .A4(new_n291_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n300_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n298_), .A2(new_n299_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n292_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(new_n299_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n292_), .A2(new_n307_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n300_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G120gat), .B(G148gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(G176gat), .B(G204gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n306_), .A2(new_n311_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT13), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(KEYINPUT13), .A3(new_n320_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G15gat), .B(G22gat), .ZN(new_n326_));
  INV_X1    g125(.A(G1gat), .ZN(new_n327_));
  INV_X1    g126(.A(G8gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT14), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G8gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(new_n291_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G231gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT17), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G127gat), .B(G155gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT16), .ZN(new_n338_));
  XOR2_X1   g137(.A(G183gat), .B(G211gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n335_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(KEYINPUT17), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n335_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT37), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n278_), .B(new_n344_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n284_), .A2(new_n325_), .A3(new_n343_), .A4(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n346_), .A2(KEYINPUT80), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(KEYINPUT80), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350_));
  INV_X1    g149(.A(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT30), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT87), .ZN(new_n355_));
  AND3_X1   g154(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G169gat), .ZN(new_n359_));
  INV_X1    g158(.A(G176gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(KEYINPUT24), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G183gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT25), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G183gat), .ZN(new_n366_));
  INV_X1    g165(.A(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT26), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT26), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G190gat), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n364_), .A2(new_n366_), .A3(new_n368_), .A4(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n361_), .A2(KEYINPUT24), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(KEYINPUT84), .A3(new_n373_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n362_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n359_), .A2(KEYINPUT22), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G169gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n379_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n379_), .B1(new_n381_), .B2(G169gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n360_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n372_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n358_), .B2(new_n389_), .ZN(new_n390_));
  NOR4_X1   g189(.A1(new_n356_), .A2(new_n357_), .A3(new_n388_), .A4(KEYINPUT86), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n386_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n355_), .B1(new_n378_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n362_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n377_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT84), .B1(new_n371_), .B2(new_n373_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n390_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n391_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n380_), .A2(new_n382_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n360_), .B(new_n384_), .C1(new_n400_), .C2(new_n379_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .A4(new_n372_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(new_n402_), .A3(KEYINPUT87), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT88), .B(G15gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n393_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n393_), .B2(new_n403_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n354_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(new_n353_), .A3(new_n408_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(KEYINPUT90), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT91), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G127gat), .B(G134gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G120gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n416_), .A2(new_n417_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT89), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT31), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n415_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT91), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n411_), .A2(new_n413_), .A3(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n415_), .A2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n349_), .B(new_n423_), .C1(new_n426_), .C2(new_n422_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n415_), .A2(new_n422_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n422_), .B1(new_n415_), .B2(new_n425_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT92), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G22gat), .B(G50gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  INV_X1    g233(.A(G141gat), .ZN(new_n435_));
  INV_X1    g234(.A(G148gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT93), .B1(G141gat), .B2(G148gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  OR2_X1    g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G141gat), .A2(G148gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n439_), .A2(new_n443_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT2), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n440_), .A2(new_n442_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n446_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT28), .B1(new_n456_), .B2(KEYINPUT29), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n456_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n433_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n457_), .A3(new_n432_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G211gat), .B(G218gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(KEYINPUT94), .A2(G197gat), .ZN(new_n467_));
  INV_X1    g266(.A(G204gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT94), .A2(G197gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT21), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(G197gat), .B2(G204gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n466_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G197gat), .A2(G204gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n467_), .A2(new_n469_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(G204gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n473_), .B1(KEYINPUT21), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n465_), .A2(new_n471_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(KEYINPUT95), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT95), .B1(new_n476_), .B2(new_n478_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n456_), .A2(KEYINPUT29), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(G78gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(new_n221_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n483_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n464_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n464_), .A2(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n460_), .A2(new_n462_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT96), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G225gat), .A2(G233gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT99), .Z(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n456_), .A2(new_n420_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n446_), .B(new_n455_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT4), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n456_), .A2(new_n420_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n499_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G29gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT100), .B(G85gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT0), .B(G57gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n498_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n512_));
  OR3_X1    g311(.A1(new_n505_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n496_), .A2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G8gat), .B(G36gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G64gat), .B(G92gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G226gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT19), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n378_), .A2(new_n392_), .A3(new_n355_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT87), .B1(new_n397_), .B2(new_n402_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n482_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n529_));
  INV_X1    g328(.A(new_n481_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n476_), .A2(KEYINPUT21), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n530_), .A2(new_n479_), .B1(new_n531_), .B2(new_n473_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n372_), .A2(KEYINPUT97), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n372_), .A2(KEYINPUT97), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n400_), .A2(new_n360_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n358_), .A2(new_n389_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n362_), .B2(new_n374_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n529_), .B1(new_n532_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n525_), .B1(new_n528_), .B2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n393_), .A2(new_n403_), .A3(new_n532_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n529_), .B1(new_n482_), .B2(new_n538_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n542_), .A2(new_n525_), .A3(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n522_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n524_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n522_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n528_), .A2(new_n525_), .A3(new_n540_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n545_), .A2(KEYINPUT27), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT102), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n532_), .B1(new_n393_), .B2(new_n403_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT20), .B1(new_n482_), .B2(new_n538_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n553_), .A2(new_n524_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n525_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n522_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n550_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT27), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n552_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI211_X1 g359(.A(KEYINPUT102), .B(KEYINPUT27), .C1(new_n557_), .C2(new_n550_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n517_), .B(new_n551_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT103), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT101), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n514_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n502_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n500_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n568_), .A2(new_n510_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n514_), .A2(new_n565_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n557_), .A2(new_n550_), .A3(new_n566_), .A4(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n548_), .A2(KEYINPUT32), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n547_), .A2(new_n549_), .A3(new_n572_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n515_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n496_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n564_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  AOI211_X1 g378(.A(KEYINPUT101), .B(new_n496_), .C1(new_n571_), .C2(new_n576_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n555_), .A2(new_n556_), .A3(new_n522_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n548_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n559_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT102), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n558_), .A2(new_n552_), .A3(new_n559_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT103), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n551_), .A4(new_n517_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n563_), .A2(new_n581_), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n551_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT104), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT104), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n593_), .B(new_n551_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n496_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n427_), .A2(new_n430_), .A3(new_n516_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n431_), .A2(new_n590_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n251_), .A2(new_n332_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT81), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n332_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n264_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n600_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(G113gat), .B(G141gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(G169gat), .B(G197gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n605_), .A2(new_n614_), .A3(new_n608_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n597_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n347_), .A2(new_n348_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n347_), .A2(KEYINPUT105), .A3(new_n348_), .A4(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n516_), .A2(G1gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n203_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n597_), .A2(new_n283_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n325_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n343_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n619_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n516_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n623_), .A2(new_n624_), .A3(new_n626_), .A4(new_n202_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1324gat));
  NAND2_X1  g437(.A1(new_n592_), .A2(new_n594_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(G8gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n623_), .A2(new_n624_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n623_), .A2(KEYINPUT108), .A3(new_n624_), .A4(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G8gat), .B1(new_n633_), .B2(new_n639_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT39), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n647_), .A3(KEYINPUT40), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1325gat));
  OAI21_X1  g451(.A(G15gat), .B1(new_n633_), .B2(new_n431_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT41), .Z(new_n654_));
  OR2_X1    g453(.A1(new_n431_), .A2(G15gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n625_), .B2(new_n655_), .ZN(G1326gat));
  OAI21_X1  g455(.A(G22gat), .B1(new_n633_), .B2(new_n578_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n578_), .A2(G22gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n625_), .B2(new_n659_), .ZN(G1327gat));
  INV_X1    g459(.A(new_n283_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n630_), .A2(new_n343_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n620_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G29gat), .B1(new_n664_), .B2(new_n515_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n345_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n267_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n282_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n344_), .B1(new_n669_), .B2(new_n278_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n666_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT43), .B1(new_n597_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n590_), .A2(new_n431_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n595_), .A2(new_n596_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n284_), .A2(new_n345_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n672_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n325_), .A2(new_n631_), .A3(new_n618_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n683_), .B(new_n680_), .C1(new_n672_), .C2(new_n678_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n515_), .A2(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n665_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688_));
  INV_X1    g487(.A(new_n639_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT109), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n639_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OR3_X1    g494(.A1(new_n663_), .A2(new_n688_), .A3(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n688_), .B1(new_n663_), .B2(new_n695_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n682_), .A2(new_n684_), .A3(new_n639_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n694_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT46), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n679_), .A2(new_n681_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n683_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n679_), .A2(KEYINPUT44), .A3(new_n681_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n689_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n698_), .B1(new_n707_), .B2(G36gat), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n708_), .A2(KEYINPUT110), .A3(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n703_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(new_n431_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n685_), .A2(G43gat), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n351_), .B1(new_n663_), .B2(new_n431_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1330gat));
  AOI21_X1  g516(.A(G50gat), .B1(new_n664_), .B2(new_n496_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n496_), .A2(G50gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n685_), .B2(new_n719_), .ZN(G1331gat));
  NAND4_X1  g519(.A1(new_n629_), .A2(new_n630_), .A3(new_n343_), .A4(new_n619_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n516_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n597_), .A2(new_n618_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(new_n630_), .A3(new_n343_), .A4(new_n671_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n516_), .A2(G57gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(G1332gat));
  INV_X1    g525(.A(new_n693_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G64gat), .B1(new_n721_), .B2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n727_), .A2(G64gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n724_), .B2(new_n731_), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n721_), .B2(new_n431_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT49), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n431_), .A2(G71gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n724_), .B2(new_n735_), .ZN(G1334gat));
  OAI21_X1  g535(.A(G78gat), .B1(new_n721_), .B2(new_n578_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT50), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n578_), .A2(G78gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n724_), .B2(new_n739_), .ZN(G1335gat));
  NOR3_X1   g539(.A1(new_n661_), .A2(new_n325_), .A3(new_n343_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n723_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n235_), .B1(new_n742_), .B2(new_n516_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT113), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n630_), .A2(new_n631_), .A3(new_n619_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n672_), .B2(new_n678_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n235_), .A3(new_n516_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n744_), .A2(new_n748_), .ZN(G1336gat));
  NAND2_X1  g548(.A1(new_n236_), .A2(new_n237_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n750_), .A3(new_n693_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n742_), .A2(new_n639_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(G92gat), .B2(new_n752_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT114), .Z(G1337gat));
  AOI21_X1  g553(.A(new_n220_), .B1(new_n746_), .B2(new_n712_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n712_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n742_), .A2(new_n756_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n755_), .A2(KEYINPUT51), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT51), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n755_), .A2(new_n761_), .A3(new_n757_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n764_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n766_), .A2(new_n759_), .A3(KEYINPUT51), .A4(new_n762_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1338gat));
  NAND4_X1  g567(.A1(new_n723_), .A2(new_n221_), .A3(new_n496_), .A4(new_n741_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n578_), .B(new_n745_), .C1(new_n672_), .C2(new_n678_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n221_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n746_), .B2(new_n496_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n770_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n745_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n679_), .A2(new_n772_), .A3(new_n496_), .A4(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G106gat), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n779_), .A2(new_n774_), .A3(KEYINPUT52), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n769_), .B1(new_n776_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT53), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n783_), .B(new_n769_), .C1(new_n776_), .C2(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1339gat));
  AOI21_X1  g584(.A(new_n299_), .B1(new_n298_), .B2(new_n305_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n306_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n298_), .A2(new_n305_), .A3(KEYINPUT55), .A4(new_n299_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n790_), .C2(new_n319_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n319_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n618_), .A2(new_n320_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n600_), .A2(new_n607_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n615_), .B1(new_n798_), .B2(new_n604_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n603_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n799_), .A2(new_n800_), .B1(new_n606_), .B2(new_n802_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n801_), .A2(new_n803_), .B1(new_n615_), .B2(new_n609_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n321_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n283_), .B1(new_n797_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT120), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  AOI211_X1 g609(.A(KEYINPUT56), .B(new_n319_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n804_), .A2(new_n320_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n793_), .A2(new_n792_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n814_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT58), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n817_), .A3(new_n677_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n809_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n806_), .A2(new_n808_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n631_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OR3_X1    g620(.A1(new_n346_), .A2(KEYINPUT54), .A3(new_n618_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT54), .B1(new_n346_), .B2(new_n618_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n516_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n595_), .A2(new_n712_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829_), .B2(new_n618_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n825_), .A2(KEYINPUT59), .A3(new_n827_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n618_), .A2(G113gat), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT121), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n830_), .B1(new_n834_), .B2(new_n836_), .ZN(G1340gat));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n325_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n829_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n325_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n838_), .ZN(G1341gat));
  INV_X1    g641(.A(G127gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n829_), .A2(new_n843_), .A3(new_n343_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n631_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n843_), .ZN(G1342gat));
  AOI21_X1  g645(.A(G134gat), .B1(new_n829_), .B2(new_n283_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT122), .B(G134gat), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n671_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n847_), .B1(new_n834_), .B2(new_n849_), .ZN(G1343gat));
  NOR3_X1   g649(.A1(new_n693_), .A2(new_n578_), .A3(new_n712_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n825_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n619_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n435_), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n325_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n436_), .ZN(G1345gat));
  NAND2_X1  g655(.A1(new_n821_), .A2(new_n824_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(new_n343_), .A3(new_n515_), .A4(new_n851_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n825_), .A2(KEYINPUT123), .A3(new_n343_), .A4(new_n851_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n852_), .B2(new_n671_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n661_), .A2(G162gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n852_), .B2(new_n867_), .ZN(G1347gat));
  NAND3_X1  g667(.A1(new_n693_), .A2(new_n578_), .A3(new_n596_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n816_), .A2(KEYINPUT58), .B1(new_n284_), .B2(new_n345_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n815_), .A2(new_n871_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n806_), .A2(new_n808_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n343_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n822_), .A2(new_n823_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n618_), .B(new_n870_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n869_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n400_), .A3(new_n618_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT62), .B1(new_n876_), .B2(G169gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT124), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(G169gat), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n879_), .A4(new_n877_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n887_), .ZN(G1348gat));
  NAND2_X1  g687(.A1(new_n878_), .A2(new_n630_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n360_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT125), .B(G176gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n889_), .B2(new_n892_), .ZN(G1349gat));
  NAND2_X1  g692(.A1(new_n878_), .A2(new_n343_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n363_), .B2(new_n894_), .ZN(G1350gat));
  NAND4_X1  g695(.A1(new_n878_), .A2(new_n283_), .A3(new_n368_), .A4(new_n370_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n878_), .A2(new_n677_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n367_), .ZN(G1351gat));
  NAND2_X1  g698(.A1(new_n431_), .A2(new_n517_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT126), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n857_), .A2(new_n693_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n618_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g704(.A1(new_n902_), .A2(new_n325_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1353gat));
  NOR2_X1   g707(.A1(new_n902_), .A2(new_n631_), .ZN(new_n909_));
  OR2_X1    g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT63), .B(G211gat), .Z(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n909_), .B2(new_n912_), .ZN(G1354gat));
  OR3_X1    g712(.A1(new_n902_), .A2(G218gat), .A3(new_n661_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G218gat), .B1(new_n902_), .B2(new_n671_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1355gat));
endmodule


