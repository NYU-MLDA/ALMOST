//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT22), .B(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT23), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT80), .ZN(new_n212_));
  OR3_X1    g011(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n210_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n208_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(new_n211_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n216_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G197gat), .B(G204gat), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT21), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT21), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n228_), .A2(KEYINPUT90), .A3(new_n229_), .A4(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n233_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT20), .B1(new_n226_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n214_), .A2(new_n223_), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n206_), .B(KEYINPUT81), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n224_), .A2(new_n215_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n207_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n239_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(KEYINPUT91), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT91), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n245_), .B(new_n233_), .C1(new_n234_), .C2(new_n236_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n203_), .B1(new_n238_), .B2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G8gat), .B(G36gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(G64gat), .B(G92gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n203_), .B1(new_n226_), .B2(new_n237_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n244_), .A2(new_n243_), .A3(new_n246_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(KEYINPUT20), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n248_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT27), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT102), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT101), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n223_), .A2(new_n224_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n214_), .A2(new_n215_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n261_), .B(new_n262_), .C1(new_n263_), .C2(new_n208_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n237_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n237_), .A2(new_n265_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT101), .B1(new_n216_), .B2(new_n225_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .A4(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(KEYINPUT20), .A3(new_n255_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n203_), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n238_), .A2(new_n247_), .A3(new_n203_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n260_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n203_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n255_), .A2(KEYINPUT20), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n276_), .B2(new_n269_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(KEYINPUT102), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n259_), .B(KEYINPUT103), .C1(new_n279_), .C2(new_n253_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT103), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT102), .B1(new_n277_), .B2(new_n272_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n271_), .A2(new_n260_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n253_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n281_), .B1(new_n284_), .B2(new_n258_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n248_), .A2(new_n256_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(new_n253_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT27), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n280_), .A2(new_n285_), .A3(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n266_), .A2(new_n267_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(G155gat), .B2(G162gat), .ZN(new_n297_));
  INV_X1    g096(.A(G141gat), .ZN(new_n298_));
  INV_X1    g097(.A(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n300_), .A2(KEYINPUT3), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(KEYINPUT3), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n304_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n297_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT1), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n300_), .B(new_n302_), .C1(new_n296_), .C2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n293_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n291_), .B1(new_n292_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n311_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT86), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(KEYINPUT86), .A3(new_n311_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(KEYINPUT29), .A3(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n291_), .B(KEYINPUT89), .Z(new_n319_));
  NAND4_X1  g118(.A1(new_n318_), .A2(new_n246_), .A3(new_n244_), .A4(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n313_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT94), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n321_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n316_), .A2(new_n317_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  AOI211_X1 g127(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n316_), .C2(new_n317_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT87), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n317_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT86), .B1(new_n308_), .B2(new_n311_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n327_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT28), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT87), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G22gat), .B(G50gat), .Z(new_n338_));
  NAND3_X1  g137(.A1(new_n330_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n330_), .B2(new_n337_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT88), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n330_), .A2(new_n337_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n338_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT88), .B1(new_n346_), .B2(new_n339_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n324_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n313_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n321_), .A2(new_n322_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n346_), .A2(new_n349_), .A3(new_n350_), .A4(new_n339_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G127gat), .B(G134gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G113gat), .B(G120gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n308_), .A2(new_n311_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n357_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n353_), .A2(new_n354_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n355_), .B2(new_n362_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n316_), .A2(new_n317_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT4), .B1(new_n360_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n316_), .A2(new_n317_), .A3(new_n364_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n367_), .B1(new_n360_), .B2(new_n365_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G85gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT0), .B(G57gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n372_), .A2(new_n380_), .A3(new_n373_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G15gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n243_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(new_n364_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G43gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n387_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n383_), .A2(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n290_), .A2(new_n352_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n379_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n356_), .B(KEYINPUT96), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n370_), .B1(new_n399_), .B2(new_n369_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n371_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n367_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT98), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT98), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n404_), .B(new_n367_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT97), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n380_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n380_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT97), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n403_), .A2(new_n405_), .A3(new_n408_), .A4(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n374_), .A2(KEYINPUT33), .A3(new_n378_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n398_), .A2(new_n287_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT32), .B(new_n253_), .C1(new_n274_), .C2(new_n278_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n253_), .A2(KEYINPUT32), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(KEYINPUT99), .Z(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n248_), .A3(new_n256_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT100), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n382_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n351_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n342_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n346_), .A2(KEYINPUT88), .A3(new_n339_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n424_), .B2(new_n324_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n321_), .B(new_n323_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n383_), .B1(new_n428_), .B2(new_n421_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n290_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n394_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n396_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G29gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G43gat), .B(G50gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT15), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G15gat), .B(G22gat), .ZN(new_n437_));
  INV_X1    g236(.A(G1gat), .ZN(new_n438_));
  INV_X1    g237(.A(G8gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT14), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G1gat), .B(G8gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n435_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G229gat), .A2(G233gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n443_), .B(new_n445_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n447_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G141gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT78), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G169gat), .B(G197gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(KEYINPUT77), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n452_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT79), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n432_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G85gat), .A2(G92gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n471_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT65), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n476_));
  INV_X1    g275(.A(G99gat), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT7), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n465_), .B1(new_n475_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT68), .ZN(new_n484_));
  INV_X1    g283(.A(G92gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n485_), .A2(KEYINPUT9), .ZN(new_n486_));
  INV_X1    g285(.A(new_n464_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(new_n462_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT9), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT64), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT9), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n491_), .A3(new_n462_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT64), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n492_), .B(new_n493_), .C1(new_n465_), .C2(new_n486_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n478_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n490_), .A2(new_n494_), .A3(new_n470_), .A4(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n498_), .A2(new_n470_), .A3(new_n472_), .A4(new_n474_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT8), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT68), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n499_), .A2(KEYINPUT67), .A3(new_n465_), .A4(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n484_), .A2(new_n497_), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G71gat), .B(G78gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT11), .ZN(new_n506_));
  XOR2_X1   g305(.A(G71gat), .B(G78gat), .Z(new_n507_));
  INV_X1    g306(.A(G64gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(G57gat), .ZN(new_n509_));
  INV_X1    g308(.A(G57gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(G64gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n511_), .A3(KEYINPUT11), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n506_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT69), .ZN(new_n516_));
  OAI211_X1 g315(.A(KEYINPUT67), .B(new_n465_), .C1(new_n475_), .C2(new_n482_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n500_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n503_), .A2(KEYINPUT70), .A3(new_n516_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT70), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n518_), .A2(new_n484_), .A3(new_n502_), .A4(new_n497_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n515_), .B(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n520_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n523_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n519_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G230gat), .ZN(new_n527_));
  INV_X1    g326(.A(G233gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n515_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n525_), .A2(new_n531_), .B1(new_n521_), .B2(new_n533_), .ZN(new_n534_));
  OAI22_X1  g333(.A1(new_n521_), .A2(new_n523_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G120gat), .B(G148gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(G176gat), .B(G204gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n538_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT13), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT13), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G190gat), .B(G218gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT74), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT36), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n503_), .A2(KEYINPUT73), .A3(new_n435_), .A4(new_n518_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n521_), .B2(new_n445_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n521_), .A2(new_n436_), .B1(new_n566_), .B2(new_n565_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n561_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n561_), .B2(new_n569_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n557_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n561_), .A2(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n567_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT36), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n556_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n561_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n572_), .A2(KEYINPUT75), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(KEYINPUT37), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n572_), .B(new_n579_), .C1(KEYINPUT75), .C2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT16), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT17), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n443_), .B(new_n591_), .Z(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n516_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n516_), .B2(new_n592_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n589_), .A2(KEYINPUT17), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT76), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n592_), .B(new_n515_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n552_), .A2(new_n585_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n461_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n382_), .A2(new_n438_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT104), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT38), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n580_), .B(KEYINPUT105), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n432_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n459_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n552_), .A2(new_n609_), .A3(new_n599_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n611_), .B2(new_n383_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n604_), .A2(KEYINPUT38), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n605_), .A2(new_n612_), .A3(new_n613_), .ZN(G1324gat));
  INV_X1    g413(.A(new_n601_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n439_), .A3(new_n290_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n352_), .A2(new_n290_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n431_), .A2(new_n382_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n290_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n382_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n620_), .A2(new_n621_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n619_), .B1(new_n622_), .B2(new_n394_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n623_), .A2(new_n290_), .A3(new_n606_), .A4(new_n610_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G8gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT106), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT106), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n628_), .A3(G8gat), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n626_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n627_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n616_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT40), .B(new_n616_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n611_), .B2(new_n431_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT41), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n601_), .A2(G15gat), .A3(new_n431_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1326gat));
  XNOR2_X1  g439(.A(new_n425_), .B(KEYINPUT107), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n608_), .A2(new_n610_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G22gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT42), .ZN(new_n644_));
  INV_X1    g443(.A(G22gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n615_), .A2(new_n645_), .A3(new_n641_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(KEYINPUT109), .ZN(new_n648_));
  INV_X1    g447(.A(new_n599_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n552_), .A2(new_n649_), .A3(new_n580_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n461_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n460_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n623_), .A2(new_n652_), .A3(new_n650_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT109), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G29gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n382_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n585_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT43), .B1(new_n432_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n623_), .A2(new_n660_), .A3(new_n585_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n552_), .A2(new_n609_), .A3(new_n649_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n662_), .A2(KEYINPUT44), .A3(new_n663_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n382_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(G29gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n668_), .B2(G29gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n657_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT44), .B1(new_n662_), .B2(new_n663_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n663_), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n665_), .B(new_n676_), .C1(new_n659_), .C2(new_n661_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n678_), .B2(new_n290_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n620_), .A2(G36gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n651_), .A2(new_n654_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n673_), .B1(new_n679_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n681_), .B(KEYINPUT45), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n675_), .A2(new_n677_), .A3(new_n620_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n685_), .B(KEYINPUT46), .C1(new_n686_), .C2(new_n674_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1329gat));
  NAND3_X1  g487(.A1(new_n651_), .A2(new_n394_), .A3(new_n654_), .ZN(new_n689_));
  INV_X1    g488(.A(G43gat), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n431_), .A2(new_n690_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n678_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n666_), .A2(new_n667_), .A3(new_n692_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT47), .B1(new_n696_), .B2(new_n691_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1330gat));
  AOI21_X1  g497(.A(G50gat), .B1(new_n655_), .B2(new_n641_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n352_), .A2(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n678_), .B2(new_n700_), .ZN(G1331gat));
  INV_X1    g500(.A(new_n552_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n702_), .A2(new_n652_), .A3(new_n599_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n608_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n383_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n585_), .A2(new_n599_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n702_), .A2(new_n459_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n623_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n510_), .A3(new_n382_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(G1332gat));
  OAI21_X1  g509(.A(G64gat), .B1(new_n704_), .B2(new_n620_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n508_), .A3(new_n290_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n704_), .B2(new_n431_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n431_), .A2(G71gat), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT110), .Z(new_n718_));
  NAND2_X1  g517(.A1(new_n708_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1334gat));
  NAND3_X1  g519(.A1(new_n608_), .A2(new_n641_), .A3(new_n703_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G78gat), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT50), .ZN(new_n723_));
  INV_X1    g522(.A(G78gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n708_), .A2(new_n724_), .A3(new_n641_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1335gat));
  NAND3_X1  g525(.A1(new_n552_), .A2(new_n609_), .A3(new_n599_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n383_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n580_), .A2(new_n649_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n623_), .A2(new_n731_), .A3(new_n707_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n732_), .A2(G85gat), .A3(new_n383_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1336gat));
  OAI21_X1  g533(.A(G92gat), .B1(new_n729_), .B2(new_n620_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n732_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n485_), .A3(new_n290_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1337gat));
  NOR2_X1   g537(.A1(new_n729_), .A2(new_n431_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n477_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n394_), .A2(new_n495_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n732_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT51), .B1(new_n740_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744_));
  OAI221_X1 g543(.A(new_n744_), .B1(new_n732_), .B2(new_n741_), .C1(new_n739_), .C2(new_n477_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1338gat));
  NAND3_X1  g545(.A1(new_n736_), .A2(new_n478_), .A3(new_n352_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n728_), .A2(new_n352_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G106gat), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT52), .B(new_n478_), .C1(new_n728_), .C2(new_n352_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(new_n747_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  INV_X1    g555(.A(KEYINPUT120), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n706_), .A2(new_n460_), .A3(new_n702_), .ZN(new_n758_));
  XOR2_X1   g557(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT54), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n600_), .A2(new_n460_), .A3(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n444_), .A2(new_n446_), .A3(new_n450_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n449_), .A2(new_n447_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n456_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT115), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n767_), .A2(KEYINPUT115), .ZN(new_n770_));
  OAI22_X1  g569(.A1(new_n769_), .A2(new_n770_), .B1(new_n456_), .B2(new_n452_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n548_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n525_), .A2(new_n531_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n521_), .A2(new_n533_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n774_), .A2(new_n524_), .A3(new_n519_), .A4(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n529_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n534_), .A2(new_n536_), .A3(KEYINPUT55), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780_));
  INV_X1    g579(.A(new_n775_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT12), .B1(new_n521_), .B2(new_n523_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n781_), .A2(new_n535_), .A3(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n784_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n537_), .A2(KEYINPUT113), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n779_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n544_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n788_), .A2(new_n789_), .A3(new_n792_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(KEYINPUT55), .A2(new_n783_), .B1(new_n776_), .B2(new_n529_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT113), .B1(new_n537_), .B2(new_n786_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n780_), .B(new_n784_), .C1(new_n534_), .C2(new_n536_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n546_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT114), .B1(new_n797_), .B2(new_n791_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n793_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n547_), .A2(new_n609_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n773_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT57), .B1(new_n803_), .B2(new_n580_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n790_), .B1(new_n788_), .B2(new_n544_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n789_), .B1(new_n788_), .B2(new_n792_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n785_), .A2(new_n787_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n792_), .B1(new_n807_), .B2(new_n794_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT114), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n772_), .B1(new_n810_), .B2(new_n801_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n580_), .A2(KEYINPUT57), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n771_), .A2(new_n547_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT58), .B(new_n813_), .C1(new_n798_), .C2(new_n808_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n585_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n811_), .A2(new_n812_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n599_), .B1(new_n804_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT119), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n599_), .C1(new_n804_), .C2(new_n819_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n764_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  NOR4_X1   g623(.A1(new_n352_), .A2(new_n290_), .A3(new_n383_), .A4(new_n431_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT117), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n757_), .B1(new_n824_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n764_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n823_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  INV_X1    g631(.A(new_n580_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n811_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n812_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n798_), .A2(new_n799_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n802_), .B1(new_n836_), .B2(new_n809_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n837_), .B2(new_n772_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n817_), .A2(new_n585_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n814_), .A2(new_n815_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n834_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n822_), .B1(new_n842_), .B2(new_n599_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n830_), .B1(new_n831_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n828_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(KEYINPUT120), .A3(new_n845_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n803_), .A2(new_n835_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n649_), .B1(new_n847_), .B2(new_n834_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n826_), .B1(new_n848_), .B2(new_n764_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT59), .ZN(new_n850_));
  INV_X1    g649(.A(G113gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n460_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n829_), .A2(new_n846_), .A3(new_n850_), .A4(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n826_), .B(new_n459_), .C1(new_n764_), .C2(new_n848_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n854_), .A2(KEYINPUT118), .A3(new_n851_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT118), .B1(new_n854_), .B2(new_n851_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n853_), .A2(KEYINPUT121), .A3(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1340gat));
  NAND3_X1  g661(.A1(new_n829_), .A2(new_n846_), .A3(new_n850_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G120gat), .B1(new_n863_), .B2(new_n702_), .ZN(new_n864_));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n702_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(KEYINPUT60), .B2(new_n865_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n849_), .B2(new_n867_), .ZN(G1341gat));
  INV_X1    g667(.A(G127gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n599_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n829_), .A2(new_n846_), .A3(new_n850_), .A4(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n849_), .B2(new_n599_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT122), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(new_n875_), .A3(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1342gat));
  OAI21_X1  g676(.A(G134gat), .B1(new_n863_), .B2(new_n658_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n606_), .A2(G134gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n849_), .B2(new_n879_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n848_), .A2(new_n764_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n620_), .A2(new_n352_), .A3(new_n382_), .A4(new_n431_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886_), .B2(new_n609_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n298_), .B(new_n459_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1344gat));
  OAI21_X1  g688(.A(G148gat), .B1(new_n886_), .B2(new_n702_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n299_), .B(new_n552_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1345gat));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(new_n886_), .B2(new_n599_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n893_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n649_), .B(new_n895_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n886_), .B2(new_n658_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n606_), .A2(G162gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1347gat));
  NAND2_X1  g700(.A1(new_n290_), .A2(new_n618_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n641_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n844_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n844_), .A2(KEYINPUT124), .A3(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(new_n204_), .A3(new_n459_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G169gat), .B1(new_n904_), .B2(new_n609_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n910_), .A2(KEYINPUT62), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(KEYINPUT62), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n909_), .B1(new_n911_), .B2(new_n912_), .ZN(G1348gat));
  NAND2_X1  g712(.A1(new_n908_), .A2(new_n552_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n881_), .A2(new_n352_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n902_), .A2(new_n205_), .A3(new_n702_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n205_), .B1(new_n915_), .B2(new_n916_), .ZN(G1349gat));
  NAND3_X1  g716(.A1(new_n290_), .A2(new_n618_), .A3(new_n649_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G183gat), .B1(new_n915_), .B2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n599_), .A2(new_n217_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n908_), .B2(new_n921_), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n908_), .A2(new_n218_), .A3(new_n607_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n658_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n210_), .B2(new_n924_), .ZN(G1351gat));
  NAND3_X1  g724(.A1(new_n621_), .A2(new_n290_), .A3(new_n431_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n881_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n459_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n552_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n931_));
  XOR2_X1   g730(.A(new_n930_), .B(new_n931_), .Z(G1353gat));
  AOI21_X1  g731(.A(new_n599_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n927_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT126), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n938_));
  XOR2_X1   g737(.A(new_n937_), .B(KEYINPUT127), .Z(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n934_), .B2(new_n939_), .ZN(G1354gat));
  INV_X1    g739(.A(G218gat), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n927_), .A2(new_n941_), .A3(new_n607_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n881_), .A2(new_n658_), .A3(new_n926_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n941_), .ZN(G1355gat));
endmodule


