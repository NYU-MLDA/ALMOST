//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_, new_n981_;
  XOR2_X1   g000(.A(G71gat), .B(G99gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT31), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT82), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  INV_X1    g005(.A(G134gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G127gat), .ZN(new_n208_));
  INV_X1    g007(.A(G127gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G134gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT81), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n206_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n209_), .A2(G134gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n207_), .A2(G127gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT81), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G113gat), .B(G120gat), .Z(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n205_), .B1(new_n214_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n212_), .A2(new_n213_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT82), .B1(new_n222_), .B2(new_n219_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n204_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G227gat), .A2(G233gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n226_), .B(G15gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT30), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n225_), .A2(new_n228_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT25), .B(G183gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT23), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(KEYINPUT24), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n233_), .A2(new_n235_), .A3(new_n239_), .A4(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n236_), .A2(KEYINPUT22), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT22), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G169gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n245_), .B2(G169gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n237_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT79), .B(new_n240_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT80), .ZN(new_n251_));
  OR2_X1    g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n235_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(G183gat), .B2(G190gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT80), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(new_n253_), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT22), .B(G169gat), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n237_), .B(new_n248_), .C1(new_n259_), .C2(new_n243_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT79), .B1(new_n260_), .B2(new_n240_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n242_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT83), .ZN(new_n263_));
  OR3_X1    g062(.A1(new_n229_), .A2(new_n230_), .A3(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G29gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT93), .B(G85gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT0), .B(G57gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n273_));
  AND3_X1   g072(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT1), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT84), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280_));
  NAND3_X1  g079(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n276_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G141gat), .B(G148gat), .Z(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288_));
  INV_X1    g087(.A(G141gat), .ZN(new_n289_));
  INV_X1    g088(.A(G148gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n291_), .A2(new_n294_), .A3(new_n295_), .A4(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n283_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n297_), .A2(KEYINPUT85), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT85), .B1(new_n297_), .B2(new_n298_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n287_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n212_), .A2(new_n213_), .A3(new_n206_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n219_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT82), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n222_), .A2(new_n219_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n205_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  OAI221_X1 g106(.A(new_n287_), .B1(new_n302_), .B2(new_n303_), .C1(new_n300_), .C2(new_n299_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n273_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT4), .B1(new_n224_), .B2(new_n301_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n308_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n311_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n272_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT33), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(KEYINPUT33), .B(new_n272_), .C1(new_n312_), .C2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n311_), .B1(new_n313_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(new_n321_), .B2(new_n313_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n311_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n271_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT91), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n234_), .A2(KEYINPUT23), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n234_), .A2(KEYINPUT23), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n326_), .B(new_n252_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT91), .B1(new_n255_), .B2(new_n256_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n240_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n259_), .B2(new_n237_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT21), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT86), .ZN(new_n335_));
  OR2_X1    g134(.A1(G197gat), .A2(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G197gat), .A2(G204gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G211gat), .B(G218gat), .Z(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G211gat), .B(G218gat), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n341_), .A2(new_n336_), .A3(new_n337_), .A4(new_n335_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n334_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n333_), .A2(new_n345_), .A3(new_n242_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT19), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT92), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n354_), .A2(new_n341_), .B1(new_n334_), .B2(new_n343_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(KEYINPUT87), .A3(new_n340_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT87), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n345_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n262_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n353_), .B1(new_n262_), .B2(new_n359_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n352_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT18), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  NAND2_X1  g165(.A1(new_n333_), .A2(new_n242_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n345_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n349_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n262_), .B2(new_n359_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n348_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n366_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n262_), .A2(new_n359_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT92), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n262_), .A2(new_n359_), .A3(new_n353_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n351_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n370_), .A2(new_n348_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n373_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n325_), .A2(new_n372_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n362_), .A2(new_n381_), .A3(new_n371_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n312_), .A2(new_n315_), .A3(new_n272_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n313_), .A2(KEYINPUT4), .ZN(new_n384_));
  INV_X1    g183(.A(new_n311_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n310_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n271_), .B1(new_n387_), .B2(new_n314_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n382_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT95), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n367_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n333_), .A2(KEYINPUT95), .A3(new_n242_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n345_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n361_), .B2(new_n360_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n368_), .B1(new_n367_), .B2(new_n390_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n349_), .B1(new_n396_), .B2(new_n392_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT96), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n348_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n370_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n348_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n381_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n320_), .A2(new_n380_), .B1(new_n389_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G228gat), .ZN(new_n405_));
  INV_X1    g204(.A(G233gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT87), .B1(new_n355_), .B2(new_n340_), .ZN(new_n409_));
  AND4_X1   g208(.A1(KEYINPUT87), .A2(new_n340_), .A3(new_n344_), .A4(new_n342_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n297_), .A2(new_n298_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n297_), .A2(new_n298_), .A3(KEYINPUT85), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n412_), .B1(new_n417_), .B2(new_n287_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n411_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n415_), .A2(new_n416_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n301_), .A2(KEYINPUT89), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n368_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n419_), .B1(new_n426_), .B2(new_n407_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT90), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n421_), .A2(new_n412_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G22gat), .B(G50gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT28), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n431_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n427_), .A2(new_n429_), .ZN(new_n436_));
  AOI211_X1 g235(.A(new_n428_), .B(new_n419_), .C1(new_n426_), .C2(new_n407_), .ZN(new_n437_));
  OAI22_X1  g236(.A1(new_n430_), .A2(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n426_), .A2(new_n407_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n428_), .B1(new_n439_), .B2(new_n419_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n427_), .A2(new_n429_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT90), .A4(new_n434_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n404_), .A2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n438_), .A2(new_n442_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT27), .B1(new_n379_), .B2(new_n372_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n375_), .A2(new_n376_), .B1(new_n397_), .B2(KEYINPUT96), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n393_), .A2(KEYINPUT20), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT96), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n401_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n402_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n373_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n372_), .A2(KEYINPUT27), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n446_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n387_), .A2(new_n271_), .A3(new_n314_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n316_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n316_), .B2(new_n457_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n445_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n266_), .B1(new_n444_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n456_), .A2(new_n443_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n266_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G8gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT74), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT72), .B(G15gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G22gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G1gat), .A2(G8gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(KEYINPUT14), .B2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n471_), .A2(new_n475_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G29gat), .B(G36gat), .Z(new_n478_));
  XOR2_X1   g277(.A(G43gat), .B(G50gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OR3_X1    g280(.A1(new_n476_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n471_), .B(new_n475_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n480_), .B(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n482_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n483_), .B(new_n480_), .ZN(new_n490_));
  OAI211_X1 g289(.A(KEYINPUT76), .B(new_n489_), .C1(new_n490_), .C2(new_n488_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n489_), .A2(KEYINPUT76), .ZN(new_n492_));
  XOR2_X1   g291(.A(G113gat), .B(G141gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT77), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G169gat), .B(G197gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n467_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT13), .ZN(new_n502_));
  INV_X1    g301(.A(G85gat), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT6), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n513_));
  INV_X1    g312(.A(G99gat), .ZN(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n507_), .B1(new_n512_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT8), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n509_), .A2(new_n511_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n517_), .A3(new_n516_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT8), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n507_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n506_), .A2(KEYINPUT9), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n527_));
  OR2_X1    g326(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n515_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n505_), .A2(KEYINPUT9), .A3(new_n506_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  XOR2_X1   g335(.A(G71gat), .B(G78gat), .Z(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n537_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n534_), .A2(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(KEYINPUT12), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT12), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n522_), .A2(new_n523_), .A3(new_n507_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n523_), .B1(new_n522_), .B2(new_n507_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n530_), .A2(new_n531_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n506_), .A2(KEYINPUT9), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n521_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT65), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n527_), .A2(new_n554_), .A3(new_n530_), .A4(new_n531_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n546_), .B1(new_n549_), .B2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n553_), .A2(new_n555_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(new_n525_), .A3(KEYINPUT66), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n545_), .B(new_n541_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT64), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n544_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n542_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(new_n543_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G120gat), .B(G148gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G176gat), .B(G204gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n566_), .A2(new_n572_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n502_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(KEYINPUT13), .A3(new_n573_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n541_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n483_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n582_), .A2(new_n583_), .A3(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(KEYINPUT17), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n582_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n549_), .A2(new_n546_), .A3(new_n556_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT66), .B1(new_n558_), .B2(new_n525_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n486_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT34), .ZN(new_n598_));
  OAI22_X1  g397(.A1(new_n533_), .A2(new_n481_), .B1(KEYINPUT35), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT68), .ZN(new_n601_));
  INV_X1    g400(.A(new_n598_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n596_), .A2(new_n600_), .A3(new_n601_), .A4(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT69), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT36), .B1(new_n609_), .B2(new_n610_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT70), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n604_), .A2(new_n601_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT68), .B1(new_n602_), .B2(new_n603_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n485_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n619_), .B(new_n620_), .C1(new_n621_), .C2(new_n599_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n605_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n613_), .B1(new_n605_), .B2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT37), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n605_), .A2(new_n622_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n613_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n622_), .A2(new_n605_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n625_), .A2(new_n631_), .A3(KEYINPUT71), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT71), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n633_), .B(KEYINPUT37), .C1(new_n623_), .C2(new_n624_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n579_), .A2(new_n593_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n501_), .A2(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT98), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT98), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n461_), .A2(G1gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(KEYINPUT38), .A3(new_n642_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n579_), .A2(new_n593_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n628_), .A2(new_n630_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n501_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n461_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n646_), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT99), .ZN(G1324gat));
  OAI21_X1  g451(.A(G8gat), .B1(new_n649_), .B2(new_n456_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n654_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n456_), .A2(G8gat), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n655_), .B(new_n656_), .C1(new_n640_), .C2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g458(.A(new_n266_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n640_), .A2(G15gat), .A3(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT101), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(KEYINPUT101), .ZN(new_n663_));
  OAI21_X1  g462(.A(G15gat), .B1(new_n649_), .B2(new_n660_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  NAND3_X1  g464(.A1(new_n662_), .A2(new_n663_), .A3(new_n665_), .ZN(G1326gat));
  OR2_X1    g465(.A1(new_n649_), .A2(new_n443_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G22gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G22gat), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n443_), .A2(G22gat), .ZN(new_n671_));
  OAI22_X1  g470(.A1(new_n669_), .A2(new_n670_), .B1(new_n640_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT102), .Z(G1327gat));
  INV_X1    g472(.A(new_n500_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(new_n576_), .A3(new_n578_), .A4(new_n593_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n467_), .A2(new_n675_), .A3(new_n648_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n461_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n675_), .B(KEYINPUT103), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n635_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n316_), .A2(new_n457_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT97), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n316_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n684_), .A2(new_n438_), .A3(new_n442_), .A4(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n366_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n377_), .A2(new_n378_), .A3(new_n373_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n366_), .B1(new_n362_), .B2(new_n371_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n687_), .A2(new_n454_), .B1(new_n690_), .B2(KEYINPUT27), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n686_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n690_), .A2(new_n325_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n375_), .A2(new_n376_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n450_), .A2(new_n694_), .A3(new_n394_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n452_), .B1(new_n695_), .B2(new_n348_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n683_), .B(new_n382_), .C1(new_n696_), .C2(new_n381_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n693_), .A2(new_n697_), .B1(new_n442_), .B2(new_n438_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n660_), .B1(new_n692_), .B2(new_n698_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n464_), .A2(new_n465_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n682_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n699_), .A2(KEYINPUT105), .A3(new_n700_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n681_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n635_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n467_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n708_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n701_), .A2(KEYINPUT106), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n679_), .B1(new_n705_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT44), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n675_), .B(new_n716_), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n706_), .B(new_n708_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT106), .B1(new_n701_), .B2(new_n710_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n702_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n635_), .A3(new_n704_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n680_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n717_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT107), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n715_), .A2(new_n725_), .B1(KEYINPUT44), .B2(new_n724_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n677_), .A2(G29gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n678_), .B1(new_n726_), .B2(new_n727_), .ZN(G1328gat));
  INV_X1    g527(.A(G36gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n726_), .B2(new_n691_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n676_), .A2(new_n729_), .A3(new_n691_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT45), .Z(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n734_), .A3(KEYINPUT46), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1329gat));
  NAND3_X1  g537(.A1(new_n726_), .A2(G43gat), .A3(new_n266_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G43gat), .B1(new_n676_), .B2(new_n266_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT108), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT47), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n741_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1330gat));
  INV_X1    g545(.A(G50gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n676_), .A2(new_n747_), .A3(new_n445_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n443_), .B1(new_n724_), .B2(KEYINPUT44), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n751_), .B1(new_n724_), .B2(KEYINPUT107), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n714_), .B(new_n717_), .C1(new_n720_), .C2(new_n723_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n749_), .B(new_n750_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G50gat), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n713_), .A2(new_n714_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n725_), .A3(new_n751_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n749_), .B1(new_n757_), .B2(new_n750_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n748_), .B1(new_n755_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT110), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n748_), .C1(new_n755_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1331gat));
  INV_X1    g562(.A(new_n579_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n467_), .A2(new_n764_), .A3(new_n674_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n592_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n635_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT111), .ZN(new_n768_));
  INV_X1    g567(.A(G57gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n677_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n648_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n766_), .A2(new_n771_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n772_), .A2(KEYINPUT112), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(KEYINPUT112), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n677_), .A3(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n770_), .B1(new_n775_), .B2(new_n769_), .ZN(G1332gat));
  INV_X1    g575(.A(G64gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n777_), .A3(new_n691_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n773_), .A2(new_n691_), .A3(new_n774_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G64gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G64gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(G1333gat));
  INV_X1    g582(.A(G71gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n768_), .A2(new_n784_), .A3(new_n266_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n773_), .A2(new_n266_), .A3(new_n774_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G71gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G71gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(G1334gat));
  INV_X1    g589(.A(G78gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n768_), .A2(new_n791_), .A3(new_n445_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n773_), .A2(new_n445_), .A3(new_n774_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(new_n794_), .A3(G78gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(G78gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(G1335gat));
  NOR3_X1   g596(.A1(new_n764_), .A2(new_n674_), .A3(new_n592_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801_), .B2(new_n461_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n765_), .A2(new_n593_), .A3(new_n771_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n677_), .A2(new_n503_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT113), .Z(G1336gat));
  OAI21_X1  g605(.A(G92gat), .B1(new_n801_), .B2(new_n456_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n691_), .A2(new_n504_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT114), .ZN(G1337gat));
  NAND3_X1  g609(.A1(new_n266_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n803_), .A2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT115), .ZN(new_n813_));
  OAI21_X1  g612(.A(G99gat), .B1(new_n801_), .B2(new_n660_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g615(.A(new_n798_), .B(new_n445_), .C1(new_n705_), .C2(new_n712_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT116), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n800_), .A2(new_n819_), .A3(new_n445_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n820_), .A3(G106gat), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT52), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n818_), .A2(new_n820_), .A3(new_n823_), .A4(G106gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n803_), .A2(G106gat), .A3(new_n443_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT53), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(new_n829_), .A3(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1339gat));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n636_), .A2(new_n500_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n563_), .A2(KEYINPUT117), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n544_), .A2(new_n560_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n836_), .A2(KEYINPUT55), .B1(new_n562_), .B2(new_n837_), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n563_), .A2(KEYINPUT117), .A3(KEYINPUT55), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n571_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT56), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n572_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n490_), .B1(G229gat), .B2(G233gat), .ZN(new_n846_));
  AND4_X1   g645(.A1(G229gat), .A2(new_n482_), .A3(G233gat), .A4(new_n487_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n496_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n574_), .A2(new_n849_), .A3(new_n499_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n842_), .A2(new_n845_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n842_), .A2(new_n845_), .A3(KEYINPUT58), .A4(new_n850_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n635_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n853_), .A2(KEYINPUT119), .A3(new_n854_), .A4(new_n635_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n849_), .A2(new_n499_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n573_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n841_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n843_), .A2(new_n864_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n862_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n859_), .B1(new_n868_), .B2(new_n771_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n868_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT57), .A3(new_n648_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n857_), .A2(new_n858_), .A3(new_n869_), .A4(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n835_), .B1(new_n872_), .B2(new_n593_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n464_), .A2(new_n660_), .A3(new_n461_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n873_), .A2(new_n500_), .A3(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n832_), .B1(new_n876_), .B2(G113gat), .ZN(new_n877_));
  INV_X1    g676(.A(G113gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n872_), .A2(new_n593_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n835_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n874_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT120), .B(new_n878_), .C1(new_n882_), .C2(new_n500_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n871_), .A2(new_n869_), .A3(new_n855_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n593_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n880_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n875_), .A2(KEYINPUT59), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n882_), .A2(KEYINPUT59), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n500_), .A2(new_n878_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n877_), .A2(new_n883_), .B1(new_n888_), .B2(new_n889_), .ZN(G1340gat));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n887_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n873_), .A2(new_n875_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G120gat), .B1(new_n894_), .B2(new_n764_), .ZN(new_n895_));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n764_), .B2(KEYINPUT60), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n892_), .B(new_n897_), .C1(KEYINPUT60), .C2(new_n896_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(new_n898_), .ZN(G1341gat));
  AOI21_X1  g698(.A(G127gat), .B1(new_n892_), .B2(new_n592_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n592_), .A2(G127gat), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n901_), .B(KEYINPUT121), .Z(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n888_), .B2(new_n902_), .ZN(G1342gat));
  OAI21_X1  g702(.A(G134gat), .B1(new_n894_), .B2(new_n682_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n892_), .A2(new_n207_), .A3(new_n771_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1343gat));
  NOR4_X1   g705(.A1(new_n691_), .A2(new_n461_), .A3(new_n443_), .A4(new_n266_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n881_), .A2(new_n674_), .A3(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g708(.A1(new_n881_), .A2(new_n579_), .A3(new_n907_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g710(.A1(new_n881_), .A2(new_n592_), .A3(new_n907_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT61), .B(G155gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1346gat));
  INV_X1    g713(.A(G162gat), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n881_), .A2(new_n915_), .A3(new_n771_), .A4(new_n907_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n881_), .A2(new_n635_), .A3(new_n907_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n915_), .ZN(G1347gat));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n835_), .B1(new_n884_), .B2(new_n593_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n691_), .A2(new_n461_), .A3(new_n266_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT122), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n443_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n920_), .A2(new_n500_), .A3(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G169gat), .B1(new_n924_), .B2(KEYINPUT123), .ZN(new_n925_));
  INV_X1    g724(.A(new_n923_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n886_), .A2(new_n674_), .A3(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n919_), .B1(new_n925_), .B2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n236_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n924_), .A2(KEYINPUT123), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n931_), .A2(KEYINPUT62), .A3(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n924_), .A2(new_n259_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(new_n933_), .A3(new_n934_), .ZN(G1348gat));
  NAND2_X1  g734(.A1(new_n881_), .A2(new_n443_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n922_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n937_), .A2(new_n237_), .A3(new_n764_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n936_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n920_), .A2(new_n923_), .ZN(new_n941_));
  AOI21_X1  g740(.A(G176gat), .B1(new_n941_), .B2(new_n579_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT124), .B1(new_n940_), .B2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n886_), .A2(new_n926_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n237_), .B1(new_n944_), .B2(new_n764_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n945_), .B(new_n946_), .C1(new_n936_), .C2(new_n939_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n943_), .A2(new_n947_), .ZN(G1349gat));
  NOR2_X1   g747(.A1(new_n873_), .A2(new_n445_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n937_), .A2(new_n593_), .ZN(new_n950_));
  AOI21_X1  g749(.A(G183gat), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n593_), .A2(new_n231_), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n941_), .A2(KEYINPUT125), .A3(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(KEYINPUT125), .B1(new_n941_), .B2(new_n952_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n951_), .A2(new_n953_), .A3(new_n954_), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n944_), .B2(new_n682_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n941_), .A2(new_n232_), .A3(new_n771_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1351gat));
  NOR2_X1   g757(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(KEYINPUT127), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n686_), .A2(new_n456_), .A3(new_n266_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n873_), .A2(new_n962_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(new_n674_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n960_), .B1(new_n964_), .B2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n965_), .ZN(new_n967_));
  INV_X1    g766(.A(new_n960_), .ZN(new_n968_));
  AOI211_X1 g767(.A(new_n967_), .B(new_n968_), .C1(new_n963_), .C2(new_n674_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n966_), .A2(new_n969_), .ZN(G1352gat));
  NAND2_X1  g769(.A1(new_n963_), .A2(new_n579_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  AND2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  OAI211_X1 g773(.A(new_n963_), .B(new_n592_), .C1(new_n973_), .C2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n963_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n976_), .A2(new_n593_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n975_), .B1(new_n977_), .B2(new_n973_), .ZN(G1354gat));
  OAI21_X1  g777(.A(G218gat), .B1(new_n976_), .B2(new_n682_), .ZN(new_n979_));
  INV_X1    g778(.A(G218gat), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n963_), .A2(new_n980_), .A3(new_n771_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n979_), .A2(new_n981_), .ZN(G1355gat));
endmodule


