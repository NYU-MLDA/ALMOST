//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_;
  INV_X1    g000(.A(KEYINPUT111), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT25), .B(G183gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT26), .B1(new_n204_), .B2(KEYINPUT82), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n203_), .B(new_n205_), .C1(new_n206_), .C2(KEYINPUT82), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT83), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT23), .ZN(new_n210_));
  OR2_X1    g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT85), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(KEYINPUT85), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n211_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT84), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n208_), .A2(new_n214_), .A3(new_n215_), .A4(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT86), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT22), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n221_), .B(G169gat), .C1(KEYINPUT87), .C2(KEYINPUT22), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT87), .A2(G169gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(new_n220_), .A3(KEYINPUT22), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT88), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n222_), .A2(new_n229_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n227_), .A2(new_n228_), .A3(new_n216_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n210_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n209_), .B2(KEYINPUT23), .ZN(new_n234_));
  OAI22_X1  g033(.A1(new_n233_), .A2(new_n234_), .B1(G183gat), .B2(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n216_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n228_), .B1(new_n238_), .B2(new_n227_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n219_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT30), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n219_), .B(KEYINPUT30), .C1(new_n239_), .C2(new_n236_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT92), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G71gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G99gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(G15gat), .B(G43gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT91), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n248_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT92), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n242_), .A2(new_n252_), .A3(new_n243_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n245_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n251_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n244_), .A2(KEYINPUT92), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT93), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G127gat), .B(G134gat), .Z(new_n258_));
  XOR2_X1   g057(.A(G113gat), .B(G120gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT31), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT95), .A2(KEYINPUT3), .ZN(new_n267_));
  INV_X1    g066(.A(G141gat), .ZN(new_n268_));
  INV_X1    g067(.A(G148gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n271_));
  OAI22_X1  g070(.A1(KEYINPUT95), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(KEYINPUT94), .A2(G141gat), .A3(G148gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT94), .B1(G141gat), .B2(G148gat), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT2), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n266_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(new_n278_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n264_), .A2(KEYINPUT1), .B1(new_n268_), .B2(new_n269_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n274_), .A2(new_n275_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n277_), .A2(KEYINPUT96), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT96), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n284_), .B(new_n266_), .C1(new_n273_), .C2(new_n276_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n260_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(new_n260_), .A3(new_n285_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT4), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G225gat), .A2(G233gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n283_), .A2(new_n285_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293_));
  INV_X1    g092(.A(new_n260_), .ZN(new_n294_));
  AND4_X1   g093(.A1(KEYINPUT104), .A2(new_n292_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT104), .B1(new_n286_), .B2(new_n293_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n289_), .B(new_n291_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n287_), .A2(new_n288_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n290_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G29gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G85gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT0), .B(G57gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n254_), .A2(KEYINPUT93), .A3(new_n256_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n261_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n263_), .B(new_n308_), .C1(new_n310_), .C2(new_n257_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT107), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT20), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT22), .B(G169gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n223_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n216_), .B(KEYINPUT101), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n317_), .A2(new_n318_), .A3(KEYINPUT102), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT102), .B1(new_n317_), .B2(new_n318_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n315_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(KEYINPUT26), .B(G190gat), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n203_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n212_), .A2(new_n217_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n324_), .B(new_n325_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT21), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT98), .B(G204gat), .ZN(new_n329_));
  INV_X1    g128(.A(G197gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n328_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G211gat), .B(G218gat), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n330_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n328_), .B1(G197gat), .B2(G204gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n331_), .A2(new_n332_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n334_), .A2(KEYINPUT21), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n333_), .A2(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n314_), .B1(new_n327_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n240_), .B2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n240_), .A2(new_n341_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT103), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n327_), .B2(new_n341_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n340_), .A2(new_n321_), .A3(new_n326_), .A4(KEYINPUT103), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n345_), .A2(new_n314_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT18), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  NAND3_X1  g156(.A1(new_n346_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT106), .ZN(new_n359_));
  INV_X1    g158(.A(new_n357_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n345_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n340_), .B(KEYINPUT99), .ZN(new_n362_));
  INV_X1    g161(.A(new_n327_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n314_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n364_), .B2(new_n347_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n343_), .A2(new_n345_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n360_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT106), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n346_), .A2(new_n353_), .A3(new_n368_), .A4(new_n357_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n359_), .A2(new_n367_), .A3(KEYINPUT27), .A4(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371_));
  INV_X1    g170(.A(new_n358_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n357_), .B1(new_n346_), .B2(new_n353_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT97), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT97), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G228gat), .ZN(new_n384_));
  INV_X1    g183(.A(G233gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n340_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n379_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n362_), .B2(new_n381_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n377_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n377_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G22gat), .B(G50gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT28), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n394_), .B(new_n396_), .Z(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n390_), .B2(KEYINPUT100), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n391_), .A2(KEYINPUT100), .A3(new_n392_), .A4(new_n397_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n313_), .B1(new_n375_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n370_), .A2(new_n374_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n404_), .A2(new_n401_), .A3(KEYINPUT107), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n312_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT32), .B(new_n357_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n357_), .A2(KEYINPUT32), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n346_), .A2(new_n353_), .A3(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n407_), .B(new_n409_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n295_), .A2(new_n296_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT105), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n289_), .A2(new_n290_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n295_), .A2(new_n296_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT105), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n304_), .B1(new_n298_), .B2(new_n291_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n373_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n358_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n297_), .A2(KEYINPUT33), .A3(new_n299_), .A4(new_n304_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n410_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n402_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n401_), .A2(new_n308_), .A3(new_n374_), .A4(new_n370_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n263_), .B1(new_n310_), .B2(new_n257_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n406_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G113gat), .B(G141gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G169gat), .B(G197gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n432_), .B(new_n433_), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT78), .B(G1gat), .Z(new_n436_));
  INV_X1    g235(.A(G8gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT14), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G1gat), .B(G8gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G29gat), .B(G36gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n446_), .A2(KEYINPUT75), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(KEYINPUT75), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G43gat), .B(G50gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n445_), .B(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G229gat), .A2(G233gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT81), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n454_), .B(KEYINPUT15), .ZN(new_n460_));
  INV_X1    g259(.A(new_n445_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n445_), .A2(new_n454_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n456_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(KEYINPUT81), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n435_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n459_), .A2(new_n466_), .A3(new_n464_), .A4(new_n434_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G230gat), .A2(G233gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G64gat), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n475_));
  XOR2_X1   g274(.A(G71gat), .B(G78gat), .Z(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n475_), .A2(new_n476_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT66), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT66), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n483_));
  AND2_X1   g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT70), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n482_), .A2(KEYINPUT6), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n480_), .A2(KEYINPUT66), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT70), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n497_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n487_), .A2(new_n494_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G85gat), .B(G92gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT8), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n505_), .A2(KEYINPUT8), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n501_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n491_), .A2(KEYINPUT67), .A3(new_n493_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n509_), .B1(new_n514_), .B2(KEYINPUT69), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT69), .ZN(new_n516_));
  AOI211_X1 g315(.A(new_n516_), .B(new_n510_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n508_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT9), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(G85gat), .A3(G92gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n520_), .B1(new_n505_), .B2(new_n519_), .ZN(new_n521_));
  OR2_X1    g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT64), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(KEYINPUT64), .A3(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT65), .B(G106gat), .Z(new_n529_));
  AOI21_X1  g328(.A(new_n521_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n512_), .A2(new_n513_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n479_), .B1(new_n518_), .B2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n533_), .A2(KEYINPUT71), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n518_), .A2(new_n479_), .A3(new_n532_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n533_), .B2(KEYINPUT71), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n472_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n532_), .A2(KEYINPUT73), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n530_), .A2(new_n531_), .A3(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n518_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n477_), .A2(KEYINPUT12), .A3(new_n478_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n532_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n485_), .A2(new_n486_), .A3(new_n511_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT67), .B1(new_n491_), .B2(new_n493_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n503_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n516_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n514_), .A2(KEYINPUT69), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n509_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n545_), .B1(new_n551_), .B2(new_n508_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n542_), .A2(new_n544_), .B1(new_n552_), .B2(new_n479_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n552_), .B2(new_n479_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n471_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n537_), .A2(KEYINPUT72), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT72), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n558_), .B(new_n472_), .C1(new_n534_), .C2(new_n536_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT13), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n564_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT74), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n567_), .A2(new_n570_), .A3(KEYINPUT74), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n431_), .A2(new_n470_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n479_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n445_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT16), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n578_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT80), .Z(new_n587_));
  INV_X1    g386(.A(KEYINPUT79), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n578_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n578_), .A2(new_n588_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT8), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n509_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n548_), .B2(new_n516_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n596_), .B2(new_n550_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n454_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n545_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT34), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT35), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n542_), .A2(new_n460_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n602_), .A2(KEYINPUT35), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n600_), .A2(new_n603_), .A3(new_n604_), .A4(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT15), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n454_), .B(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n518_), .B2(new_n541_), .ZN(new_n609_));
  OAI211_X1 g408(.A(KEYINPUT35), .B(new_n602_), .C1(new_n609_), .C2(new_n599_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT76), .ZN(new_n613_));
  XOR2_X1   g412(.A(G134gat), .B(G162gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n606_), .A2(new_n616_), .A3(new_n610_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(KEYINPUT77), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(KEYINPUT37), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT37), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n619_), .B(new_n620_), .C1(KEYINPUT77), .C2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n592_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OR3_X1    g426(.A1(new_n575_), .A2(KEYINPUT108), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n308_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT108), .B1(new_n575_), .B2(new_n627_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n628_), .A2(new_n436_), .A3(new_n629_), .A4(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n573_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n574_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n470_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n592_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n621_), .B(KEYINPUT110), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n431_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n308_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n202_), .B1(new_n635_), .B2(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n631_), .A2(new_n633_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(KEYINPUT111), .A3(new_n634_), .A4(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1324gat));
  NAND3_X1  g449(.A1(new_n639_), .A2(new_n643_), .A3(new_n404_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G8gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n654_), .A3(G8gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n628_), .A2(new_n437_), .A3(new_n404_), .A4(new_n630_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1325gat));
  NOR2_X1   g460(.A1(new_n644_), .A2(new_n429_), .ZN(new_n662_));
  INV_X1    g461(.A(G15gat), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n662_), .A2(KEYINPUT113), .A3(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT113), .B1(new_n662_), .B2(new_n663_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n575_), .A2(new_n627_), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT93), .B(new_n261_), .C1(new_n254_), .C2(new_n256_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n310_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n257_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n663_), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n664_), .A2(KEYINPUT41), .A3(new_n665_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n668_), .A2(new_n674_), .A3(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n644_), .B2(new_n402_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n669_), .A2(new_n679_), .A3(new_n401_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1327gat));
  NOR2_X1   g480(.A1(new_n640_), .A2(new_n621_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n575_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n629_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n623_), .A2(new_n625_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n375_), .A2(new_n402_), .A3(new_n313_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT107), .B1(new_n404_), .B2(new_n401_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n311_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n673_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n686_), .B(new_n688_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT114), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n431_), .A2(KEYINPUT114), .A3(new_n686_), .A4(new_n688_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT43), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n696_), .A3(new_n698_), .ZN(new_n699_));
  NOR4_X1   g498(.A1(new_n636_), .A2(new_n637_), .A3(new_n640_), .A4(new_n638_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT44), .B1(new_n699_), .B2(new_n700_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n629_), .A2(G29gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n685_), .B1(new_n703_), .B2(new_n704_), .ZN(G1328gat));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n684_), .A2(new_n706_), .A3(new_n404_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT45), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n701_), .A2(new_n702_), .A3(new_n375_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n706_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n708_), .B(KEYINPUT46), .C1(new_n709_), .C2(new_n706_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  NAND2_X1  g513(.A1(new_n673_), .A2(G43gat), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n701_), .A2(new_n702_), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G43gat), .B1(new_n684_), .B2(new_n673_), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n716_), .A2(KEYINPUT47), .A3(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT47), .B1(new_n716_), .B2(new_n717_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1330gat));
  AOI21_X1  g519(.A(G50gat), .B1(new_n684_), .B2(new_n401_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n401_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n703_), .B2(new_n722_), .ZN(G1331gat));
  NOR2_X1   g522(.A1(new_n636_), .A2(new_n637_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n470_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n643_), .ZN(new_n726_));
  INV_X1    g525(.A(G57gat), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n308_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n431_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n627_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT115), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT115), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n629_), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n728_), .B1(new_n733_), .B2(new_n727_), .ZN(G1332gat));
  INV_X1    g533(.A(G64gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(new_n735_), .A3(new_n404_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737_));
  INV_X1    g536(.A(new_n726_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n404_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n739_), .B2(G64gat), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT48), .B(new_n735_), .C1(new_n738_), .C2(new_n404_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n740_), .B2(new_n741_), .ZN(G1333gat));
  OAI21_X1  g541(.A(G71gat), .B1(new_n726_), .B2(new_n429_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT49), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT49), .ZN(new_n745_));
  INV_X1    g544(.A(new_n730_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n429_), .A2(G71gat), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n744_), .A2(new_n745_), .B1(new_n746_), .B2(new_n747_), .ZN(G1334gat));
  INV_X1    g547(.A(G78gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n730_), .A2(new_n749_), .A3(new_n401_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n738_), .A2(new_n401_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G78gat), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT50), .B(new_n749_), .C1(new_n738_), .C2(new_n401_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(G1335gat));
  AOI211_X1 g554(.A(new_n640_), .B(new_n470_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n699_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n308_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n729_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n682_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n308_), .A2(G85gat), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT116), .ZN(G1336gat));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n404_), .A3(new_n682_), .ZN(new_n765_));
  INV_X1    g564(.A(G92gat), .ZN(new_n766_));
  INV_X1    g565(.A(new_n757_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n404_), .A2(G92gat), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT117), .Z(new_n769_));
  AOI22_X1  g568(.A1(new_n765_), .A2(new_n766_), .B1(new_n767_), .B2(new_n769_), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n757_), .B2(new_n429_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n673_), .A2(new_n528_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n760_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(KEYINPUT118), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n773_), .B(new_n775_), .ZN(G1338gat));
  NAND4_X1  g575(.A1(new_n759_), .A2(new_n529_), .A3(new_n401_), .A4(new_n682_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n699_), .A2(new_n401_), .A3(new_n756_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G106gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G106gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n777_), .B(new_n784_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  AOI21_X1  g585(.A(new_n470_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(new_n626_), .A3(new_n788_), .ZN(new_n789_));
  OR2_X1    g588(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n787_), .A2(new_n626_), .B1(new_n790_), .B2(new_n788_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n621_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n638_), .A2(new_n566_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  INV_X1    g597(.A(new_n563_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n471_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n556_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n553_), .A2(KEYINPUT55), .A3(new_n471_), .A4(new_n555_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n798_), .B(new_n799_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n538_), .A2(new_n540_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n544_), .B1(new_n597_), .B2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n535_), .C1(new_n533_), .C2(KEYINPUT12), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n801_), .B1(new_n807_), .B2(new_n472_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n472_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n803_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n563_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n798_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n804_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT120), .A3(new_n798_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n797_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n462_), .A2(new_n818_), .A3(new_n463_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n456_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n434_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n469_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n568_), .B2(new_n564_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n795_), .B1(new_n817_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n814_), .B1(new_n827_), .B2(KEYINPUT56), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(KEYINPUT56), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n816_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n825_), .B1(new_n830_), .B2(new_n796_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n794_), .B1(new_n831_), .B2(new_n793_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n557_), .A2(new_n559_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n824_), .B1(new_n833_), .B2(new_n799_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n802_), .A2(new_n803_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT56), .B1(new_n835_), .B2(new_n563_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n836_), .B2(new_n804_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT58), .B(new_n834_), .C1(new_n836_), .C2(new_n804_), .ZN(new_n840_));
  AND4_X1   g639(.A1(KEYINPUT122), .A2(new_n839_), .A3(new_n688_), .A4(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n687_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT122), .B1(new_n842_), .B2(new_n840_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n826_), .B(new_n832_), .C1(new_n841_), .C2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n792_), .B1(new_n844_), .B2(new_n592_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n403_), .A2(new_n405_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n673_), .A2(new_n629_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n845_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n842_), .A2(new_n840_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n832_), .A2(new_n826_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n592_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n792_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n848_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT123), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n792_), .B1(new_n852_), .B2(new_n592_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n857_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n850_), .B1(new_n859_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G113gat), .B1(new_n863_), .B2(new_n638_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n845_), .A2(new_n849_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n470_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1340gat));
  XOR2_X1   g667(.A(KEYINPUT124), .B(G120gat), .Z(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n863_), .B2(new_n724_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n724_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n865_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1341gat));
  OAI21_X1  g673(.A(G127gat), .B1(new_n863_), .B2(new_n592_), .ZN(new_n875_));
  INV_X1    g674(.A(G127gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n865_), .A2(new_n876_), .A3(new_n640_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1342gat));
  OAI21_X1  g677(.A(G134gat), .B1(new_n863_), .B2(new_n687_), .ZN(new_n879_));
  INV_X1    g678(.A(G134gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n641_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n865_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1343gat));
  NOR2_X1   g682(.A1(new_n841_), .A2(new_n843_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n832_), .A2(new_n826_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n592_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n854_), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n673_), .A2(new_n308_), .A3(new_n402_), .A4(new_n404_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT125), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  INV_X1    g689(.A(new_n888_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n845_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n470_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G141gat), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n268_), .B(new_n470_), .C1(new_n889_), .C2(new_n892_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1344gat));
  INV_X1    g695(.A(new_n724_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G148gat), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n269_), .B(new_n897_), .C1(new_n889_), .C2(new_n892_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1345gat));
  OAI21_X1  g700(.A(new_n640_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n903_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n640_), .B(new_n905_), .C1(new_n889_), .C2(new_n892_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1346gat));
  INV_X1    g706(.A(G162gat), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n908_), .B(new_n881_), .C1(new_n889_), .C2(new_n892_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n887_), .A2(KEYINPUT125), .A3(new_n888_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n890_), .B1(new_n845_), .B2(new_n891_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n687_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n909_), .B1(new_n908_), .B2(new_n912_), .ZN(G1347gat));
  NOR3_X1   g712(.A1(new_n311_), .A2(new_n401_), .A3(new_n375_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n638_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G169gat), .B1(new_n860_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n831_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n919_), .A2(new_n795_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n640_), .B1(new_n920_), .B2(new_n832_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n316_), .B(new_n916_), .C1(new_n921_), .C2(new_n792_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n918_), .A2(new_n922_), .A3(KEYINPUT62), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n924_), .B(G169gat), .C1(new_n860_), .C2(new_n917_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT126), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n923_), .A2(new_n928_), .A3(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1348gat));
  NOR2_X1   g729(.A1(new_n860_), .A2(new_n915_), .ZN(new_n931_));
  AOI21_X1  g730(.A(G176gat), .B1(new_n931_), .B2(new_n897_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n845_), .A2(new_n915_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n724_), .A2(new_n223_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1349gat));
  AOI21_X1  g734(.A(G183gat), .B1(new_n933_), .B2(new_n640_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n592_), .A2(new_n203_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n931_), .B2(new_n937_), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n931_), .A2(new_n323_), .A3(new_n881_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n860_), .A2(new_n687_), .A3(new_n915_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n204_), .B2(new_n940_), .ZN(G1351gat));
  NAND3_X1  g740(.A1(new_n404_), .A2(new_n308_), .A3(new_n401_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n845_), .A2(new_n673_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n470_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g744(.A(G204gat), .B1(new_n943_), .B2(new_n897_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n329_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n943_), .A2(new_n897_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n946_), .B1(new_n947_), .B2(new_n948_), .ZN(G1353gat));
  AOI21_X1  g748(.A(new_n592_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n943_), .A2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT127), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n951_), .B(new_n954_), .ZN(G1354gat));
  INV_X1    g754(.A(G218gat), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n943_), .A2(new_n956_), .A3(new_n881_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n943_), .A2(new_n688_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n956_), .ZN(G1355gat));
endmodule


