//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(G204gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G197gat), .ZN(new_n203_));
  INV_X1    g002(.A(G197gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G204gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT21), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n206_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT97), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n208_), .B(new_n207_), .C1(new_n210_), .C2(new_n212_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT25), .B(G183gat), .Z(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT26), .ZN(new_n219_));
  AND2_X1   g018(.A1(KEYINPUT88), .A2(G190gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT88), .A2(G190gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT26), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT89), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT89), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n224_), .B(KEYINPUT26), .C1(new_n220_), .C2(new_n221_), .ZN(new_n225_));
  AOI211_X1 g024(.A(new_n217_), .B(new_n219_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  INV_X1    g026(.A(G176gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT24), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT90), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT23), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n223_), .A2(new_n225_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n217_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n219_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT90), .ZN(new_n242_));
  INV_X1    g041(.A(new_n231_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n232_), .A2(new_n237_), .A3(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n227_), .A2(new_n228_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G169gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(new_n228_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(KEYINPUT91), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n220_), .A2(new_n221_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n234_), .B1(new_n251_), .B2(G183gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(KEYINPUT91), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n216_), .B1(new_n245_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT20), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n239_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n229_), .B(KEYINPUT101), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n234_), .A2(KEYINPUT102), .A3(new_n236_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT102), .B1(new_n234_), .B2(new_n236_), .ZN(new_n261_));
  OAI221_X1 g060(.A(new_n258_), .B1(new_n259_), .B2(new_n230_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n248_), .B(KEYINPUT103), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n234_), .B1(G183gat), .B2(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n216_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n255_), .A2(new_n256_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT106), .B1(new_n269_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n245_), .A2(new_n254_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n267_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n268_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT20), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT106), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n271_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n245_), .A2(new_n254_), .A3(new_n216_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n256_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n272_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n273_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT18), .B(G64gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G92gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT32), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n283_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G225gat), .A2(G233gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  AND2_X1   g093(.A1(KEYINPUT96), .A2(KEYINPUT2), .ZN(new_n295_));
  NOR2_X1   g094(.A1(KEYINPUT96), .A2(KEYINPUT2), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(G141gat), .B(G148gat), .C1(KEYINPUT96), .C2(KEYINPUT2), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .A4(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n308_), .A3(new_n305_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n300_), .A2(KEYINPUT95), .ZN(new_n310_));
  NAND3_X1  g109(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n311_), .A2(new_n294_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n300_), .A2(KEYINPUT95), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n307_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G120gat), .ZN(new_n316_));
  OR2_X1    g115(.A1(G127gat), .A2(G134gat), .ZN(new_n317_));
  INV_X1    g116(.A(G113gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G127gat), .A2(G134gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n316_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G113gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(G120gat), .A3(new_n320_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n315_), .A2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n307_), .A2(new_n323_), .A3(new_n314_), .A4(new_n326_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(KEYINPUT105), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT105), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n315_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n293_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n328_), .A2(KEYINPUT4), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n292_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n330_), .A2(new_n291_), .A3(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G85gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(G1gat), .B(G29gat), .Z(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n337_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n280_), .A2(new_n281_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n271_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT104), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n269_), .A2(new_n272_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n272_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT104), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .A4(new_n288_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n290_), .A2(new_n343_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n287_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT33), .B1(new_n337_), .B2(new_n342_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357_));
  AOI211_X1 g156(.A(new_n357_), .B(new_n341_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .A4(new_n287_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n333_), .A2(new_n292_), .A3(new_n334_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n291_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n361_), .A2(new_n342_), .A3(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n355_), .A2(new_n359_), .A3(new_n360_), .A4(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n352_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT30), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n245_), .A2(new_n366_), .A3(new_n254_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n245_), .B2(new_n254_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n327_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n274_), .A2(KEYINPUT30), .ZN(new_n370_));
  INV_X1    g169(.A(new_n327_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n245_), .A2(new_n366_), .A3(new_n254_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G15gat), .B(G43gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n369_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G71gat), .B(G99gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT94), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n381_), .B(new_n383_), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n376_), .A2(new_n377_), .A3(new_n385_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n367_), .A2(new_n368_), .A3(new_n327_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n371_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n374_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n369_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n384_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G78gat), .B(G106gat), .Z(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT98), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n395_), .A2(new_n267_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n307_), .B2(new_n314_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n397_), .B(KEYINPUT98), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n400_), .A2(new_n216_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n394_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n401_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n395_), .A2(new_n267_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n397_), .A2(new_n396_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(new_n400_), .B2(new_n216_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n393_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT100), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT99), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n403_), .A2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G22gat), .B(G50gat), .Z(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT28), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n416_), .A2(new_n309_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n417_), .B2(new_n399_), .ZN(new_n418_));
  AND4_X1   g217(.A1(new_n415_), .A2(new_n307_), .A3(new_n399_), .A4(new_n314_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n414_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT28), .B1(new_n315_), .B2(KEYINPUT29), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n415_), .A3(new_n399_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n413_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n410_), .B1(new_n412_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n405_), .A2(new_n407_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT99), .B1(new_n427_), .B2(new_n394_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n428_), .A2(KEYINPUT100), .A3(new_n424_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n409_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n412_), .A2(new_n410_), .A3(new_n425_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT100), .B1(new_n428_), .B2(new_n424_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n403_), .A4(new_n408_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n365_), .A2(new_n392_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n355_), .A2(new_n360_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n283_), .A2(new_n354_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(KEYINPUT27), .A3(new_n360_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n385_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(new_n433_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n389_), .A2(new_n384_), .A3(new_n390_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n442_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n438_), .B(new_n440_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n435_), .B1(new_n446_), .B2(new_n343_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G57gat), .B(G64gat), .Z(new_n448_));
  INV_X1    g247(.A(KEYINPUT11), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n449_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G71gat), .A2(G78gat), .ZN(new_n452_));
  INV_X1    g251(.A(G71gat), .ZN(new_n453_));
  INV_X1    g252(.A(G78gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT69), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT69), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n451_), .A2(new_n458_), .A3(new_n452_), .A4(new_n455_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n450_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n457_), .A2(new_n459_), .A3(new_n450_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G99gat), .ZN(new_n464_));
  INV_X1    g263(.A(G106gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT66), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(G99gat), .B2(G106gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT67), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G99gat), .A2(G106gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT67), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n466_), .A2(new_n468_), .A3(new_n478_), .A4(new_n469_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G85gat), .A2(G92gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n480_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n474_), .A2(new_n475_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(KEYINPUT9), .B2(new_n484_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT65), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT10), .B(G99gat), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(G106gat), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n481_), .A2(KEYINPUT9), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n490_), .A2(new_n491_), .A3(new_n493_), .A4(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G85gat), .ZN(new_n496_));
  INV_X1    g295(.A(G92gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(KEYINPUT9), .A3(new_n481_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n499_), .A2(new_n494_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n492_), .A2(G106gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT65), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n495_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n487_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n480_), .A2(new_n484_), .A3(new_n504_), .A4(new_n485_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n488_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n463_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G230gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT64), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT70), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n463_), .A2(new_n506_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT12), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n463_), .A2(KEYINPUT12), .A3(new_n506_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT70), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(new_n509_), .C1(new_n463_), .C2(new_n506_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n511_), .A2(new_n514_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n507_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n512_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n510_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G120gat), .B(G148gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT73), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT74), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G176gat), .B(G204gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n525_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n522_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n518_), .A2(new_n521_), .A3(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT13), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(KEYINPUT13), .A3(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(G8gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT81), .B(G22gat), .ZN(new_n541_));
  INV_X1    g340(.A(G15gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT82), .B(G1gat), .Z(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT14), .B1(new_n544_), .B2(new_n540_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G1gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n546_), .A2(G1gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n540_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(G8gat), .A3(new_n547_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT76), .B(G43gat), .ZN(new_n554_));
  INV_X1    g353(.A(G50gat), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G29gat), .B(G36gat), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n555_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n553_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n564_));
  OAI211_X1 g363(.A(G229gat), .B(G233gat), .C1(new_n562_), .C2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n561_), .B(KEYINPUT15), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n566_), .B(new_n567_), .C1(new_n569_), .C2(new_n553_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n227_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(new_n204_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n565_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n539_), .A2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n447_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n462_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(new_n460_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n461_), .A2(new_n462_), .A3(new_n581_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n552_), .A4(new_n550_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n584_), .A2(new_n585_), .B1(new_n552_), .B2(new_n550_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT83), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G127gat), .B(G155gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n594_), .A2(KEYINPUT17), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n584_), .A2(new_n585_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n553_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT83), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n586_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n589_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT85), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n589_), .A2(KEYINPUT85), .A3(new_n595_), .A4(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n597_), .A2(KEYINPUT86), .A3(new_n586_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT86), .B1(new_n597_), .B2(new_n586_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n594_), .B(KEYINPUT17), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n604_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT87), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT87), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n611_), .A3(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT75), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT34), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT35), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n568_), .A2(new_n506_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n488_), .A2(new_n503_), .A3(new_n561_), .A4(new_n505_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(KEYINPUT77), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(KEYINPUT77), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n618_), .B(new_n619_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n616_), .A2(new_n617_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n620_), .B(KEYINPUT77), .ZN(new_n626_));
  INV_X1    g425(.A(new_n624_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n618_), .A4(new_n619_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT80), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(G134gat), .ZN(new_n632_));
  INV_X1    g431(.A(G162gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT36), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT80), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n625_), .A2(new_n636_), .A3(new_n628_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n634_), .A2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT78), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n625_), .A2(new_n628_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT37), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT79), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n642_), .B(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n629_), .B2(new_n635_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n643_), .A2(new_n644_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n613_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n580_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n343_), .A3(new_n544_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT38), .ZN(new_n652_));
  INV_X1    g451(.A(new_n609_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n447_), .A2(new_n643_), .A3(new_n579_), .A4(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n343_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n656_), .ZN(G1324gat));
  NAND2_X1  g456(.A1(new_n438_), .A2(new_n440_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G8gat), .B1(new_n654_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n661_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(KEYINPUT39), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n650_), .A2(new_n540_), .A3(new_n658_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n660_), .A2(new_n661_), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT108), .B(KEYINPUT109), .Z(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT40), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n668_), .B(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n654_), .B2(new_n392_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT110), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n672_), .A2(KEYINPUT110), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n392_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n650_), .A2(new_n542_), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n679_), .A3(new_n680_), .ZN(G1326gat));
  OAI21_X1  g480(.A(G22gat), .B1(new_n654_), .B2(new_n434_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT42), .ZN(new_n683_));
  INV_X1    g482(.A(G22gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n650_), .A2(new_n684_), .A3(new_n442_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(G29gat), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n613_), .A2(new_n578_), .A3(new_n539_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n434_), .B1(new_n386_), .B2(new_n391_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(new_n655_), .A3(new_n438_), .A4(new_n440_), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT43), .B(new_n648_), .C1(new_n692_), .C2(new_n435_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  INV_X1    g493(.A(new_n648_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n447_), .B2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n688_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT44), .B(new_n688_), .C1(new_n693_), .C2(new_n696_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n687_), .B1(new_n701_), .B2(new_n343_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n613_), .A2(new_n643_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n580_), .A2(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n704_), .A2(G29gat), .A3(new_n655_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n702_), .A2(new_n705_), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n699_), .A2(new_n658_), .A3(new_n700_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n699_), .A2(KEYINPUT111), .A3(new_n658_), .A4(new_n700_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(G36gat), .A3(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n704_), .A2(G36gat), .A3(new_n659_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT45), .Z(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n711_), .A2(KEYINPUT46), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  NAND4_X1  g517(.A1(new_n699_), .A2(G43gat), .A3(new_n678_), .A4(new_n700_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n720_));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n704_), .B2(new_n392_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n720_), .B1(new_n719_), .B2(new_n722_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n719_), .A2(new_n722_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT47), .B1(new_n729_), .B2(new_n723_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n727_), .A2(new_n730_), .ZN(G1330gat));
  AOI21_X1  g530(.A(new_n555_), .B1(new_n701_), .B2(new_n442_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n704_), .A2(G50gat), .A3(new_n434_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1331gat));
  AOI21_X1  g533(.A(new_n577_), .B1(new_n692_), .B2(new_n435_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT113), .Z(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(new_n539_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n649_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G57gat), .B1(new_n739_), .B2(new_n343_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n735_), .A2(new_n643_), .A3(new_n539_), .A4(new_n613_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(new_n655_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(G57gat), .B2(new_n742_), .ZN(G1332gat));
  OAI21_X1  g542(.A(G64gat), .B1(new_n741_), .B2(new_n659_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT48), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n659_), .A2(G64gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n738_), .B2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n741_), .B2(new_n392_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT114), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT114), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(KEYINPUT49), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT49), .B1(new_n749_), .B2(new_n750_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n678_), .A2(new_n453_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT115), .ZN(new_n754_));
  OAI22_X1  g553(.A1(new_n751_), .A2(new_n752_), .B1(new_n738_), .B2(new_n754_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n741_), .B2(new_n434_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n442_), .A2(new_n454_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n738_), .B2(new_n758_), .ZN(G1335gat));
  OR2_X1    g558(.A1(new_n693_), .A2(new_n696_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n539_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n613_), .A2(new_n761_), .A3(new_n577_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n343_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G85gat), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n737_), .A2(new_n496_), .A3(new_n343_), .A4(new_n703_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(G1336gat));
  AND3_X1   g568(.A1(new_n763_), .A2(G92gat), .A3(new_n658_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n737_), .A2(new_n703_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n658_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n770_), .B1(new_n773_), .B2(new_n497_), .ZN(G1337gat));
  AOI21_X1  g573(.A(new_n464_), .B1(new_n763_), .B2(new_n678_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n392_), .A2(new_n492_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n772_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n771_), .A2(new_n492_), .A3(new_n392_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT51), .B1(new_n780_), .B2(new_n775_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1338gat));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n442_), .B(new_n762_), .C1(new_n693_), .C2(new_n696_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(G106gat), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n785_), .A3(G106gat), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n434_), .A2(G106gat), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n736_), .A2(new_n539_), .A3(new_n703_), .A4(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n784_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n786_), .A2(new_n785_), .A3(G106gat), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n784_), .B(new_n792_), .C1(new_n794_), .C2(new_n787_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n783_), .B1(new_n793_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n792_), .B1(new_n794_), .B2(new_n787_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT117), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .A3(new_n795_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n658_), .A2(new_n655_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n445_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n522_), .A2(new_n529_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n577_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n514_), .A2(new_n519_), .A3(new_n515_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n510_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n518_), .A2(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n514_), .A2(new_n515_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n812_), .A2(KEYINPUT55), .A3(new_n511_), .A4(new_n517_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n806_), .A2(KEYINPUT119), .A3(new_n510_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n809_), .A2(new_n811_), .A3(new_n813_), .A4(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n529_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n529_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n805_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n567_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n566_), .B1(new_n569_), .B2(new_n553_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n567_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n574_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n575_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n535_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n643_), .B1(new_n820_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT57), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n529_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT56), .B1(new_n815_), .B2(new_n529_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n577_), .B(new_n804_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n826_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n643_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n829_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n815_), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n529_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n825_), .A3(new_n804_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n818_), .A2(new_n819_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n839_), .B(KEYINPUT58), .C1(new_n840_), .C2(KEYINPUT120), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n830_), .A2(new_n831_), .A3(KEYINPUT120), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n838_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n844_), .A3(new_n695_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n836_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n609_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n539_), .A2(new_n577_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n649_), .A2(new_n848_), .A3(new_n849_), .A4(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n613_), .A2(new_n850_), .A3(new_n648_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT118), .B1(new_n852_), .B2(KEYINPUT54), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(KEYINPUT54), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n803_), .B1(new_n847_), .B2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n577_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n803_), .A2(KEYINPUT121), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n803_), .A2(KEYINPUT121), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n613_), .B1(new_n836_), .B2(new_n845_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n851_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n859_), .B(new_n860_), .C1(new_n861_), .C2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n858_), .A2(new_n865_), .B1(KEYINPUT122), .B2(new_n318_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  OAI21_X1  g666(.A(G113gat), .B1(new_n578_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n857_), .B1(new_n866_), .B2(new_n868_), .ZN(G1340gat));
  OAI21_X1  g668(.A(new_n316_), .B1(new_n761_), .B2(KEYINPUT60), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT123), .Z(new_n871_));
  OAI211_X1 g670(.A(new_n856_), .B(new_n871_), .C1(KEYINPUT60), .C2(new_n316_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n761_), .B1(new_n858_), .B2(new_n865_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n316_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n856_), .B2(new_n613_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT124), .B(G127gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n858_), .B2(new_n865_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n653_), .ZN(G1342gat));
  INV_X1    g677(.A(new_n643_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G134gat), .B1(new_n856_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n858_), .A2(new_n865_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n695_), .A2(G134gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT125), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n880_), .B1(new_n881_), .B2(new_n883_), .ZN(G1343gat));
  AOI21_X1  g683(.A(new_n653_), .B1(new_n836_), .B2(new_n845_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n444_), .B(new_n802_), .C1(new_n885_), .C2(new_n862_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n577_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n539_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g690(.A(new_n690_), .B1(new_n847_), .B2(new_n855_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT61), .B(G155gat), .Z(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n892_), .A2(new_n613_), .A3(new_n802_), .A4(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n613_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n893_), .B1(new_n886_), .B2(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n895_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1346gat));
  NOR3_X1   g700(.A1(new_n886_), .A2(new_n633_), .A3(new_n648_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n887_), .A2(new_n879_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n633_), .B2(new_n903_), .ZN(G1347gat));
  OR2_X1    g703(.A1(new_n861_), .A2(new_n862_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n659_), .A2(new_n343_), .A3(new_n689_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G169gat), .B1(new_n907_), .B2(new_n578_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n907_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n577_), .A3(new_n247_), .ZN(new_n912_));
  OAI211_X1 g711(.A(KEYINPUT62), .B(G169gat), .C1(new_n907_), .C2(new_n578_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n912_), .A3(new_n913_), .ZN(G1348gat));
  OAI21_X1  g713(.A(new_n228_), .B1(new_n907_), .B2(new_n761_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n659_), .A2(new_n343_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n445_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n847_), .B2(new_n855_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(G176gat), .A3(new_n539_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n915_), .A2(new_n919_), .ZN(G1349gat));
  AOI21_X1  g719(.A(G183gat), .B1(new_n918_), .B2(new_n613_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n609_), .A2(new_n239_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n911_), .B2(new_n922_), .ZN(G1350gat));
  OAI21_X1  g722(.A(G190gat), .B1(new_n907_), .B2(new_n648_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n879_), .A2(new_n257_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n907_), .B2(new_n925_), .ZN(G1351gat));
  NAND2_X1  g725(.A1(new_n892_), .A2(new_n916_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n928_), .A2(new_n204_), .A3(new_n577_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G197gat), .B1(new_n927_), .B2(new_n578_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1352gat));
  AOI21_X1  g730(.A(G204gat), .B1(new_n928_), .B2(new_n539_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n927_), .A2(new_n202_), .A3(new_n761_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1353gat));
  XOR2_X1   g733(.A(KEYINPUT63), .B(G211gat), .Z(new_n935_));
  NAND3_X1  g734(.A1(new_n928_), .A2(new_n653_), .A3(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n927_), .B2(new_n609_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1354gat));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n927_), .A2(new_n940_), .A3(new_n648_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n928_), .A2(new_n879_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1355gat));
endmodule


