//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_;
  AND2_X1   g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(KEYINPUT8), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n214_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n211_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(new_n209_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n211_), .A3(new_n221_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n217_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT10), .B(G99gat), .Z(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n206_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT9), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(G85gat), .A3(G92gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n229_), .A2(new_n230_), .A3(new_n212_), .A4(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n203_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n211_), .ZN(new_n235_));
  AND2_X1   g034(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n236_));
  NOR2_X1   g035(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n238_), .A2(new_n224_), .A3(new_n207_), .A4(new_n208_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n226_), .B1(new_n239_), .B2(new_n214_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n214_), .A2(new_n215_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n203_), .B(new_n233_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G78gat), .Z(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n234_), .A2(new_n244_), .A3(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n233_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT66), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(new_n243_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n202_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n254_), .A2(KEYINPUT12), .A3(new_n252_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n253_), .A2(new_n202_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n252_), .B1(new_n234_), .B2(new_n244_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT68), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n256_), .A2(new_n265_), .A3(KEYINPUT12), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n260_), .B(new_n261_), .C1(new_n264_), .C2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT5), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G176gat), .B(G204gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n259_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n259_), .A2(KEYINPUT69), .A3(new_n267_), .A4(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n259_), .A2(new_n267_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n271_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT13), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT14), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT79), .B(G1gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(G8gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT80), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G8gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n292_), .B(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G29gat), .B(G36gat), .Z(new_n296_));
  XOR2_X1   g095(.A(G43gat), .B(G50gat), .Z(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n292_), .B(new_n293_), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n298_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G229gat), .A2(G233gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n298_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n300_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n308_), .B2(new_n305_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G113gat), .B(G141gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G169gat), .B(G197gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n309_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G231gat), .A2(G233gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT81), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n301_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(new_n252_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G127gat), .B(G155gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT16), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G183gat), .B(G211gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT17), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT82), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT83), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n317_), .A2(new_n322_), .A3(new_n321_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n326_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n286_), .A2(new_n313_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n303_), .A2(new_n254_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n255_), .A2(new_n299_), .A3(new_n243_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G232gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT34), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n336_), .A2(KEYINPUT35), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(KEYINPUT35), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n337_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT73), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G190gat), .B(G218gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT74), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G134gat), .B(G162gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT36), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n349_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT75), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n341_), .A2(new_n343_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G169gat), .ZN(new_n362_));
  INV_X1    g161(.A(G176gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OR3_X1    g163(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT26), .B(G190gat), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT23), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n368_), .A2(new_n369_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n375_), .A2(new_n370_), .A3(G183gat), .A4(G190gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n371_), .ZN(new_n377_));
  OAI221_X1 g176(.A(new_n376_), .B1(G183gat), .B2(G190gat), .C1(new_n377_), .C2(new_n375_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G169gat), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n367_), .A2(new_n374_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n381_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G127gat), .B(G134gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G113gat), .B(G120gat), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n386_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT85), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n385_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n384_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT31), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n393_), .B(new_n398_), .Z(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT19), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT88), .B(G197gat), .ZN(new_n402_));
  INV_X1    g201(.A(G204gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT21), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(G197gat), .B2(G204gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT89), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n404_), .A2(KEYINPUT89), .A3(new_n406_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G211gat), .B(G218gat), .Z(new_n412_));
  OR2_X1    g211(.A1(G197gat), .A2(G204gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n412_), .B1(new_n414_), .B2(new_n405_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n414_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n412_), .A2(KEYINPUT21), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n411_), .A2(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n369_), .B(KEYINPUT91), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n368_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n376_), .B1(new_n377_), .B2(new_n375_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n366_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n377_), .B1(G183gat), .B2(G190gat), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n420_), .A2(new_n422_), .B1(new_n380_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT20), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n411_), .A2(new_n415_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n416_), .A2(new_n417_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n426_), .A2(new_n381_), .A3(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n401_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT92), .ZN(new_n430_));
  XOR2_X1   g229(.A(G8gat), .B(G36gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n426_), .A2(new_n427_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n381_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n401_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n418_), .A2(new_n424_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n438_), .A2(KEYINPUT20), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n442_), .B(new_n401_), .C1(new_n425_), .C2(new_n428_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n430_), .A2(new_n435_), .A3(new_n441_), .A4(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT27), .ZN(new_n445_));
  OR3_X1    g244(.A1(new_n425_), .A2(new_n428_), .A3(new_n401_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n438_), .A2(KEYINPUT20), .A3(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n401_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n435_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT100), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(KEYINPUT100), .A3(new_n450_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n445_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G22gat), .B(G50gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT86), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n459_), .B1(G155gat), .B2(G162gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G141gat), .A2(G148gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT3), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G141gat), .A2(G148gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT2), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n462_), .A2(KEYINPUT87), .A3(new_n464_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n460_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n461_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n463_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n459_), .A2(KEYINPUT1), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n473_), .B1(new_n459_), .B2(KEYINPUT1), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT29), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n477_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n457_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n481_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(new_n479_), .A3(new_n456_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(new_n484_), .A3(KEYINPUT90), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n436_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490_));
  INV_X1    g289(.A(G78gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(new_n206_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n489_), .B(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n487_), .A2(new_n488_), .A3(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G29gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G85gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT0), .B(G57gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G225gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT95), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n392_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n475_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n460_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n468_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT87), .B1(new_n462_), .B2(new_n464_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n387_), .A2(new_n388_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n501_), .B1(new_n502_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(new_n509_), .A3(KEYINPUT4), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n392_), .B(new_n513_), .C1(new_n469_), .C2(new_n475_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n501_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n499_), .B(new_n511_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n499_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n510_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n488_), .A2(new_n494_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n495_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n443_), .A2(new_n441_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n426_), .A2(new_n381_), .A3(new_n427_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(KEYINPUT20), .C1(new_n418_), .C2(new_n424_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n442_), .B1(new_n527_), .B2(new_n401_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n450_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(KEYINPUT94), .A3(new_n444_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n531_), .B(new_n450_), .C1(new_n525_), .C2(new_n528_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n530_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT102), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n530_), .A2(KEYINPUT102), .A3(new_n532_), .A4(new_n533_), .ZN(new_n537_));
  AOI211_X1 g336(.A(new_n455_), .B(new_n524_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n495_), .A2(new_n523_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n435_), .A2(KEYINPUT32), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT98), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n430_), .A2(new_n441_), .A3(new_n443_), .A4(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n449_), .A2(new_n544_), .ZN(new_n545_));
  AND4_X1   g344(.A1(KEYINPUT99), .A2(new_n521_), .A3(new_n543_), .A4(new_n545_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n517_), .A2(new_n520_), .B1(new_n449_), .B2(new_n544_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT99), .B1(new_n547_), .B2(new_n543_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n530_), .A2(new_n532_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT33), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n520_), .A2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(KEYINPUT33), .B(new_n518_), .C1(new_n519_), .C2(new_n510_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n512_), .A2(new_n516_), .A3(new_n514_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n502_), .A2(new_n509_), .A3(new_n501_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n499_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n554_), .A2(KEYINPUT97), .A3(new_n499_), .A4(new_n555_), .ZN(new_n559_));
  AND4_X1   g358(.A1(new_n552_), .A2(new_n553_), .A3(new_n558_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n550_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n540_), .B1(new_n549_), .B2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n399_), .B1(new_n538_), .B2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n455_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n399_), .A2(new_n521_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n539_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n359_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n331_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n521_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(G1gat), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n280_), .A2(new_n281_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n285_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT71), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n282_), .A2(KEYINPUT71), .A3(new_n285_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n313_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n352_), .B(KEYINPUT78), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n344_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n357_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT37), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n354_), .A2(new_n584_), .A3(new_n357_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n578_), .A2(new_n579_), .A3(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n522_), .A2(new_n288_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n592_), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT103), .B1(new_n592_), .B2(KEYINPUT38), .ZN(new_n594_));
  OAI221_X1 g393(.A(new_n570_), .B1(KEYINPUT38), .B2(new_n592_), .C1(new_n593_), .C2(new_n594_), .ZN(G1324gat));
  INV_X1    g394(.A(G8gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n564_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n331_), .A2(new_n597_), .A3(new_n567_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(G8gat), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT104), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT104), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(new_n603_), .A3(G8gat), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n601_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n602_), .B1(new_n601_), .B2(new_n604_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n598_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(KEYINPUT40), .B(new_n598_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1325gat));
  INV_X1    g410(.A(new_n399_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n395_), .B1(new_n568_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT41), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n590_), .A2(new_n395_), .A3(new_n612_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1326gat));
  INV_X1    g415(.A(G22gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n568_), .B2(new_n540_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT42), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n590_), .A2(new_n617_), .A3(new_n540_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1327gat));
  INV_X1    g420(.A(KEYINPUT107), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n521_), .A2(G29gat), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT43), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n586_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n586_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n536_), .A2(new_n537_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n455_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n524_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n547_), .A2(new_n543_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n547_), .A2(KEYINPUT99), .A3(new_n543_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n561_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n539_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n612_), .B1(new_n632_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n566_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n628_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n627_), .A2(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n286_), .A2(new_n313_), .A3(new_n587_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT44), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n625_), .A2(new_n626_), .A3(new_n624_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT43), .B1(new_n641_), .B2(KEYINPUT105), .ZN(new_n647_));
  OAI211_X1 g446(.A(KEYINPUT44), .B(new_n644_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n644_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n627_), .B2(new_n642_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n623_), .B(new_n645_), .C1(new_n650_), .C2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n330_), .A2(new_n359_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n579_), .A2(new_n573_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n521_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n622_), .B1(new_n654_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n659_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n650_), .A2(new_n653_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n645_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT107), .B(new_n661_), .C1(new_n664_), .C2(new_n623_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n660_), .A2(new_n665_), .ZN(G1328gat));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n597_), .B1(new_n652_), .B2(KEYINPUT44), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n662_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n658_), .A2(new_n668_), .A3(new_n597_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT45), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n667_), .B1(new_n671_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n669_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n676_));
  OAI211_X1 g475(.A(KEYINPUT46), .B(new_n673_), .C1(new_n676_), .C2(new_n668_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1329gat));
  NAND2_X1  g477(.A1(new_n612_), .A2(G43gat), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n679_), .B(new_n645_), .C1(new_n650_), .C2(new_n653_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G43gat), .B1(new_n658_), .B2(new_n612_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT47), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683_));
  INV_X1    g482(.A(new_n681_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n683_), .B(new_n684_), .C1(new_n664_), .C2(new_n679_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1330gat));
  AOI21_X1  g485(.A(G50gat), .B1(new_n658_), .B2(new_n540_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n664_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n540_), .A2(G50gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n688_), .B2(new_n689_), .ZN(G1331gat));
  OAI21_X1  g489(.A(new_n313_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n286_), .A3(new_n589_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(G57gat), .A3(new_n522_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n313_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n330_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT71), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n698_), .B2(new_n575_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n567_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT108), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n577_), .A2(new_n702_), .A3(new_n567_), .A4(new_n696_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n703_), .A3(new_n521_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n694_), .B1(new_n704_), .B2(G57gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT109), .ZN(G1332gat));
  OR3_X1    g505(.A1(new_n693_), .A2(G64gat), .A3(new_n564_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n701_), .A2(new_n703_), .A3(new_n597_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G64gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G64gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT110), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n707_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1333gat));
  OR3_X1    g515(.A1(new_n693_), .A2(G71gat), .A3(new_n399_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n701_), .A2(new_n703_), .A3(new_n612_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT49), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G71gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G71gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1334gat));
  NAND3_X1  g521(.A1(new_n701_), .A2(new_n703_), .A3(new_n540_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT50), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G78gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G78gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n540_), .A2(new_n491_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n725_), .A2(new_n726_), .B1(new_n693_), .B2(new_n727_), .ZN(G1335gat));
  AOI21_X1  g527(.A(new_n655_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n692_), .A3(KEYINPUT111), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n656_), .B1(new_n698_), .B2(new_n575_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n691_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G85gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n521_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n286_), .A2(new_n313_), .A3(new_n330_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n643_), .A2(KEYINPUT112), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n627_), .A2(new_n739_), .A3(new_n642_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n521_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n736_), .B1(new_n742_), .B2(new_n735_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n734_), .B2(new_n597_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n745_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n597_), .A2(G92gat), .ZN(new_n748_));
  AOI22_X1  g547(.A1(new_n746_), .A2(new_n747_), .B1(new_n741_), .B2(new_n748_), .ZN(G1337gat));
  NAND2_X1  g548(.A1(new_n612_), .A2(new_n228_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n734_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT114), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n734_), .A2(new_n754_), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n741_), .A2(new_n612_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n756_), .B(new_n757_), .C1(new_n758_), .C2(new_n205_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n757_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n754_), .B1(new_n734_), .B2(new_n751_), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT114), .B(new_n750_), .C1(new_n730_), .C2(new_n733_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n205_), .B1(new_n741_), .B2(new_n612_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n759_), .A2(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n734_), .A2(new_n206_), .A3(new_n540_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  OAI21_X1  g567(.A(G106gat), .B1(new_n768_), .B2(KEYINPUT116), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n737_), .A2(new_n539_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n643_), .B2(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n768_), .A2(KEYINPUT116), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n771_), .A2(new_n772_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n767_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT53), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n767_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1339gat));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  INV_X1    g579(.A(new_n312_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n309_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n783_));
  INV_X1    g582(.A(new_n305_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n300_), .B2(new_n307_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n785_), .B2(new_n312_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n300_), .A2(new_n304_), .A3(new_n784_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OR3_X1    g587(.A1(new_n785_), .A2(new_n783_), .A3(new_n312_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n782_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n277_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n262_), .A2(KEYINPUT68), .A3(new_n263_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n265_), .B1(new_n256_), .B2(KEYINPUT12), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n253_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n260_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n267_), .A2(KEYINPUT55), .ZN(new_n799_));
  INV_X1    g598(.A(new_n260_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n261_), .ZN(new_n803_));
  AOI221_X4 g602(.A(new_n793_), .B1(new_n798_), .B2(new_n202_), .C1(new_n799_), .C2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n799_), .A2(new_n803_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n798_), .A2(new_n202_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT118), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n792_), .B(new_n271_), .C1(new_n804_), .C2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n791_), .A2(new_n808_), .ZN(new_n809_));
  AND4_X1   g608(.A1(new_n802_), .A2(new_n796_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n802_), .B1(new_n801_), .B2(new_n261_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n793_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n805_), .A2(KEYINPUT118), .A3(new_n806_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n272_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n792_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n780_), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n271_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT56), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n808_), .A4(new_n791_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n628_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n792_), .B1(new_n815_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n313_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n280_), .A2(new_n790_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n359_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n821_), .B1(new_n828_), .B2(KEYINPUT57), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n830_), .B(new_n359_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n330_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n588_), .A2(new_n286_), .A3(new_n695_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  NOR4_X1   g635(.A1(new_n597_), .A2(new_n540_), .A3(new_n522_), .A4(new_n399_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(G113gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n695_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n838_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n836_), .A2(KEYINPUT59), .A3(new_n837_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n313_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n845_), .B2(new_n840_), .ZN(G1340gat));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n839_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n578_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n847_), .ZN(G1341gat));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n839_), .A2(new_n852_), .A3(new_n587_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n330_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n852_), .ZN(G1342gat));
  INV_X1    g654(.A(G134gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n839_), .A2(new_n856_), .A3(new_n359_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n586_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1343gat));
  NOR4_X1   g658(.A1(new_n597_), .A2(new_n539_), .A3(new_n522_), .A4(new_n612_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n836_), .A2(new_n695_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n836_), .A2(new_n577_), .A3(new_n860_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g663(.A1(new_n836_), .A2(new_n860_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n330_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT61), .B(G155gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  OAI21_X1  g667(.A(G162gat), .B1(new_n865_), .B2(new_n586_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n358_), .A2(G162gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n865_), .B2(new_n870_), .ZN(G1347gat));
  INV_X1    g670(.A(KEYINPUT22), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n597_), .A2(new_n565_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT121), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n874_), .A2(new_n695_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n836_), .A2(new_n872_), .A3(new_n539_), .A4(new_n875_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n876_), .A2(KEYINPUT62), .A3(new_n362_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(KEYINPUT62), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n836_), .A2(new_n539_), .A3(new_n875_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n362_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n877_), .B1(new_n878_), .B2(new_n881_), .ZN(G1348gat));
  AOI21_X1  g681(.A(new_n540_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n883_), .A2(new_n363_), .A3(new_n286_), .A4(new_n874_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n883_), .A2(new_n577_), .A3(new_n874_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n363_), .ZN(G1349gat));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n587_), .A3(new_n874_), .ZN(new_n887_));
  MUX2_X1   g686(.A(new_n368_), .B(G183gat), .S(new_n887_), .Z(G1350gat));
  NAND3_X1  g687(.A1(new_n883_), .A2(new_n628_), .A3(new_n874_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G190gat), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n883_), .A2(new_n419_), .A3(new_n359_), .A4(new_n874_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1351gat));
  NOR2_X1   g691(.A1(new_n524_), .A2(new_n612_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT122), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n564_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n836_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(G197gat), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n896_), .A2(new_n313_), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n695_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT123), .B(G197gat), .Z(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n901_), .B2(new_n902_), .ZN(G1352gat));
  NOR2_X1   g702(.A1(new_n896_), .A2(new_n578_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1353gat));
  AOI21_X1  g705(.A(new_n330_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n900_), .A2(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n900_), .A2(new_n907_), .A3(new_n911_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1354gat));
  INV_X1    g714(.A(G218gat), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n896_), .A2(new_n916_), .A3(new_n586_), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n836_), .A2(new_n359_), .A3(new_n895_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919_));
  AOI21_X1  g718(.A(G218gat), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT127), .B1(new_n896_), .B2(new_n358_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n917_), .B1(new_n920_), .B2(new_n921_), .ZN(G1355gat));
endmodule


