//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n204_), .B2(G106gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n203_), .A2(KEYINPUT64), .A3(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n205_), .A2(new_n211_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  OR3_X1    g016(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  XOR2_X1   g019(.A(G85gat), .B(G92gat), .Z(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n216_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n216_), .B(KEYINPUT66), .C1(new_n222_), .C2(new_n223_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G71gat), .B(G78gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n229_), .A2(new_n231_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n226_), .A2(new_n227_), .A3(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n224_), .A2(KEYINPUT12), .A3(new_n236_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n238_), .B(new_n239_), .C1(new_n240_), .C2(KEYINPUT12), .ZN(new_n241_));
  INV_X1    g040(.A(G230gat), .ZN(new_n242_));
  INV_X1    g041(.A(G233gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n240_), .A2(KEYINPUT12), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n238_), .A2(new_n239_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248_));
  INV_X1    g047(.A(new_n244_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .A4(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n238_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n244_), .B1(new_n251_), .B2(new_n240_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n245_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G120gat), .B(G148gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT5), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G176gat), .B(G204gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n245_), .A2(new_n250_), .A3(new_n252_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT13), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(KEYINPUT13), .A3(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G127gat), .B(G155gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT16), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G183gat), .B(G211gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G1gat), .B(G8gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G15gat), .ZN(new_n275_));
  INV_X1    g074(.A(G22gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G15gat), .A2(G22gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G1gat), .A2(G8gat), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n277_), .A2(new_n278_), .B1(KEYINPUT14), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n274_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G231gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n236_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n272_), .B(KEYINPUT70), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(new_n280_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(new_n282_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n237_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n271_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n284_), .A2(new_n288_), .A3(new_n270_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT17), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(KEYINPUT17), .B(new_n271_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT68), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G43gat), .B(G50gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT15), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n286_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n281_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G229gat), .A2(G233gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n300_), .A2(new_n281_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n303_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n304_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311_));
  XOR2_X1   g110(.A(G113gat), .B(G141gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT74), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G169gat), .B(G197gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n305_), .B(new_n309_), .C1(KEYINPUT73), .C2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n266_), .A2(new_n296_), .A3(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G113gat), .B(G120gat), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n322_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT79), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT75), .B(KEYINPUT23), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n329_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n328_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(KEYINPUT76), .A2(G169gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(KEYINPUT76), .A2(G169gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT22), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT77), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n341_), .B(KEYINPUT22), .C1(new_n337_), .C2(new_n338_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n343_));
  AOI21_X1  g142(.A(G176gat), .B1(new_n343_), .B2(G169gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n336_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G183gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT25), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G183gat), .ZN(new_n350_));
  INV_X1    g149(.A(G190gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT26), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT26), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G190gat), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n348_), .A2(new_n350_), .A3(new_n352_), .A4(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(KEYINPUT24), .A3(new_n327_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n355_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n331_), .A2(KEYINPUT23), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n346_), .A2(KEYINPUT30), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT30), .B1(new_n346_), .B2(new_n365_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n326_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n346_), .A2(new_n365_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n336_), .A2(new_n345_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT30), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(KEYINPUT79), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G227gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G71gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G99gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(G15gat), .B(G43gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT78), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n378_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n375_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT31), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n374_), .A2(new_n381_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n381_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n366_), .A2(new_n367_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n382_), .B1(new_n388_), .B2(KEYINPUT79), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT31), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n386_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n325_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n384_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n387_), .A2(new_n389_), .A3(KEYINPUT31), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT80), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n325_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n386_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G57gat), .B(G85gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT94), .ZN(new_n402_));
  INV_X1    g201(.A(G1gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n405_));
  INV_X1    g204(.A(G29gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n404_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n410_), .B(KEYINPUT92), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(KEYINPUT1), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT1), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n416_), .A2(KEYINPUT82), .A3(G155gat), .A4(G162gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(new_n413_), .B2(KEYINPUT1), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G141gat), .ZN(new_n421_));
  INV_X1    g220(.A(G148gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(KEYINPUT81), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(G141gat), .B2(G148gat), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n423_), .A2(new_n425_), .B1(G141gat), .B2(G148gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n420_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n413_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n428_), .A2(new_n414_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n421_), .A2(new_n422_), .A3(KEYINPUT3), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT3), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(G141gat), .B2(G148gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n430_), .A2(new_n432_), .B1(new_n433_), .B2(KEYINPUT83), .ZN(new_n434_));
  AND3_X1   g233(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT2), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n435_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n429_), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT84), .B1(new_n427_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n429_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n430_), .A2(new_n432_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n433_), .A2(KEYINPUT83), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n435_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n433_), .B2(KEYINPUT83), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n443_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n420_), .A2(new_n426_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n442_), .A2(new_n452_), .A3(new_n398_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n427_), .A2(new_n441_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n325_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n323_), .A2(KEYINPUT91), .A3(new_n324_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT4), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n453_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n412_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n453_), .A2(new_n410_), .A3(new_n458_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT95), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT95), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n453_), .A2(new_n458_), .A3(new_n466_), .A4(new_n410_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n409_), .B1(new_n463_), .B2(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n453_), .A2(new_n461_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n461_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n411_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n472_), .A2(new_n408_), .A3(new_n465_), .A4(new_n467_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n394_), .A2(new_n400_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n477_));
  INV_X1    g276(.A(G218gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G211gat), .ZN(new_n479_));
  INV_X1    g278(.A(G211gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G218gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(G197gat), .A2(G204gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G197gat), .A2(G204gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n482_), .A2(new_n485_), .A3(new_n486_), .A4(KEYINPUT21), .ZN(new_n487_));
  OR2_X1    g286(.A1(G197gat), .A2(G204gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G197gat), .A2(G204gat), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n488_), .A2(new_n486_), .A3(KEYINPUT21), .A4(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n479_), .A2(new_n481_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT21), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT85), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT85), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n497_), .B(new_n494_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n485_), .A2(KEYINPUT21), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n477_), .B1(new_n372_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT22), .B(G169gat), .ZN(new_n504_));
  INV_X1    g303(.A(G176gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n328_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(new_n363_), .B2(new_n334_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT24), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n359_), .A2(KEYINPUT88), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n327_), .B(new_n357_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n356_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n333_), .A2(new_n355_), .A3(new_n511_), .A4(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n507_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n503_), .B1(new_n515_), .B2(new_n501_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT19), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n507_), .A2(new_n514_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n483_), .A2(new_n484_), .A3(new_n494_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(KEYINPUT85), .B2(new_n495_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n522_), .A2(new_n498_), .B1(new_n492_), .B2(new_n487_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n523_), .A3(KEYINPUT89), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n502_), .A2(new_n516_), .A3(new_n519_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n520_), .A2(new_n523_), .A3(KEYINPUT89), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT89), .B1(new_n520_), .B2(new_n523_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n530_), .A2(KEYINPUT98), .A3(new_n519_), .A4(new_n502_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n501_), .A2(new_n507_), .A3(new_n514_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n533_), .B(KEYINPUT20), .C1(new_n372_), .C2(new_n501_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n534_), .B2(new_n518_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT20), .B1(new_n520_), .B2(new_n523_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n501_), .B1(new_n346_), .B2(new_n365_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n532_), .B(new_n518_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n527_), .B(new_n531_), .C1(new_n535_), .C2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G8gat), .B(G36gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G64gat), .B(G92gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT99), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n540_), .A2(KEYINPUT99), .A3(new_n546_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n502_), .A2(new_n516_), .A3(new_n524_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n518_), .ZN(new_n552_));
  OR3_X1    g351(.A1(new_n536_), .A2(new_n537_), .A3(new_n518_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n545_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT27), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n549_), .A2(new_n550_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT27), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n552_), .A2(new_n545_), .A3(new_n553_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n545_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT87), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G22gat), .B(G50gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT28), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n442_), .A2(new_n452_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n564_), .ZN(new_n568_));
  AOI211_X1 g367(.A(KEYINPUT29), .B(new_n568_), .C1(new_n442_), .C2(new_n452_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n562_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n442_), .A2(new_n452_), .A3(KEYINPUT29), .ZN(new_n571_));
  AND2_X1   g370(.A1(G228gat), .A2(G233gat), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n501_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n523_), .B1(new_n454_), .B2(new_n566_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n571_), .A2(new_n573_), .B1(new_n574_), .B2(new_n572_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G78gat), .B(G106gat), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n567_), .A2(new_n569_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n579_), .B2(KEYINPUT87), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n427_), .A2(new_n441_), .A3(KEYINPUT84), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n450_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n566_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n568_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n565_), .A2(new_n566_), .A3(new_n564_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(KEYINPUT87), .A3(new_n585_), .A4(new_n578_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n576_), .B1(new_n580_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n584_), .A2(KEYINPUT87), .A3(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n577_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n590_), .A2(new_n570_), .A3(new_n575_), .A4(new_n586_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n557_), .A2(new_n561_), .A3(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n476_), .A2(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n540_), .A2(KEYINPUT99), .A3(new_n546_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT99), .B1(new_n540_), .B2(new_n546_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n555_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n475_), .A2(new_n592_), .A3(new_n561_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT100), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n474_), .B1(new_n591_), .B2(new_n588_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n557_), .A2(new_n601_), .A3(new_n602_), .A4(new_n561_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n545_), .A2(KEYINPUT32), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n552_), .A2(new_n553_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n552_), .A2(KEYINPUT96), .A3(new_n553_), .A4(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n540_), .A2(KEYINPUT32), .A3(new_n545_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n474_), .A3(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n559_), .A2(new_n560_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n473_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n468_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n615_), .A2(KEYINPUT33), .A3(new_n408_), .A4(new_n472_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n410_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n409_), .B(new_n617_), .C1(new_n412_), .C2(new_n459_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n612_), .A2(new_n614_), .A3(new_n616_), .A4(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n611_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n593_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n600_), .A2(new_n603_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n394_), .A2(new_n400_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n595_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n301_), .A2(new_n224_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n226_), .A2(new_n227_), .A3(new_n300_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT35), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n627_), .A2(new_n628_), .B1(KEYINPUT36), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT69), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n627_), .B2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n625_), .A2(KEYINPUT69), .A3(new_n626_), .A4(new_n635_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n632_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n631_), .A2(KEYINPUT36), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n632_), .A2(new_n638_), .A3(new_n643_), .A4(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n624_), .A2(KEYINPUT103), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT103), .B1(new_n624_), .B2(new_n646_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n320_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT104), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(KEYINPUT104), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n475_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n642_), .A2(KEYINPUT37), .A3(new_n644_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n294_), .A2(KEYINPUT72), .A3(new_n295_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT72), .B1(new_n294_), .B2(new_n295_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT37), .B1(new_n642_), .B2(new_n644_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n654_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n319_), .ZN(new_n661_));
  NOR4_X1   g460(.A1(new_n624_), .A2(new_n660_), .A3(new_n661_), .A4(new_n265_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n474_), .B(KEYINPUT101), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n403_), .A3(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n653_), .A2(new_n667_), .ZN(G1324gat));
  INV_X1    g467(.A(G8gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n557_), .A2(new_n561_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n662_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n649_), .A2(new_n670_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n673_), .B2(G8gat), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT39), .B(new_n669_), .C1(new_n649_), .C2(new_n670_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1325gat));
  INV_X1    g477(.A(new_n623_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n662_), .A2(new_n275_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n681_), .B2(G15gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1326gat));
  NAND3_X1  g483(.A1(new_n662_), .A2(new_n276_), .A3(new_n592_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n592_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(G22gat), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G22gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n624_), .A2(new_n661_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n657_), .A2(new_n646_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n265_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n474_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n657_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n265_), .A2(new_n661_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n622_), .A2(new_n623_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n595_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n654_), .A2(new_n658_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n699_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n624_), .A2(KEYINPUT43), .A3(new_n703_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n698_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT106), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  INV_X1    g508(.A(new_n698_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n557_), .A2(new_n561_), .A3(new_n601_), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n711_), .A2(KEYINPUT100), .B1(new_n593_), .B2(new_n620_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n679_), .B1(new_n712_), .B2(new_n603_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n699_), .B(new_n704_), .C1(new_n713_), .C2(new_n595_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n624_), .B2(new_n703_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n710_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n708_), .A2(new_n709_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(KEYINPUT44), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n663_), .A2(new_n406_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n696_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  INV_X1    g523(.A(new_n670_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n695_), .A2(KEYINPUT45), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n728_));
  INV_X1    g527(.A(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n694_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n725_), .B1(new_n716_), .B2(KEYINPUT44), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n709_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT106), .B(new_n710_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n731_), .B1(new_n735_), .B2(G36gat), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n724_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(G36gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n719_), .B2(new_n732_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT107), .B(KEYINPUT46), .C1(new_n740_), .C2(new_n731_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1329gat));
  OAI211_X1 g541(.A(new_n679_), .B(new_n720_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G43gat), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n694_), .A2(G43gat), .A3(new_n623_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n744_), .A2(KEYINPUT47), .A3(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n695_), .B2(new_n592_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n592_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n721_), .B2(new_n752_), .ZN(G1331gat));
  NOR4_X1   g552(.A1(new_n624_), .A2(new_n660_), .A3(new_n319_), .A4(new_n266_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G57gat), .B1(new_n754_), .B2(new_n664_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n265_), .A2(new_n661_), .A3(new_n697_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT108), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT108), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT109), .B(G57gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n475_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n755_), .B1(new_n760_), .B2(new_n762_), .ZN(G1332gat));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n764_), .A3(new_n670_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n758_), .A2(new_n670_), .A3(new_n759_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G64gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G64gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(G1333gat));
  INV_X1    g569(.A(G71gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n754_), .A2(new_n771_), .A3(new_n679_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n758_), .A2(new_n679_), .A3(new_n759_), .ZN(new_n773_));
  XOR2_X1   g572(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(G71gat), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G71gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n754_), .A2(new_n778_), .A3(new_n592_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n758_), .A2(new_n592_), .A3(new_n759_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(G78gat), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G78gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(G1335gat));
  NOR4_X1   g583(.A1(new_n624_), .A2(new_n266_), .A3(new_n319_), .A4(new_n692_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G85gat), .B1(new_n785_), .B2(new_n664_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n714_), .A2(new_n715_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n265_), .A2(new_n661_), .A3(new_n657_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT112), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n475_), .A2(new_n207_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n786_), .B1(new_n791_), .B2(new_n792_), .ZN(G1336gat));
  AOI21_X1  g592(.A(G92gat), .B1(new_n785_), .B2(new_n670_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n670_), .A2(G92gat), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT113), .Z(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n791_), .B2(new_n796_), .ZN(G1337gat));
  NAND3_X1  g596(.A1(new_n785_), .A2(new_n203_), .A3(new_n679_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT114), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(new_n679_), .A3(new_n789_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(G99gat), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(G1338gat));
  NAND3_X1  g602(.A1(new_n785_), .A2(new_n214_), .A3(new_n592_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n787_), .A2(new_n592_), .A3(new_n789_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(G106gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(G106gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g609(.A1(new_n266_), .A2(new_n659_), .A3(new_n661_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n241_), .A2(new_n814_), .A3(new_n244_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n244_), .B2(new_n241_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n245_), .A2(new_n250_), .A3(new_n814_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n257_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n257_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n302_), .A2(new_n303_), .A3(new_n308_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n308_), .B1(new_n306_), .B2(new_n303_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n315_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n310_), .A2(new_n317_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n260_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n823_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n829_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n703_), .B1(new_n834_), .B2(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n319_), .A2(new_n260_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT117), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n319_), .A2(new_n840_), .A3(new_n260_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n261_), .A2(new_n828_), .ZN(new_n844_));
  OAI221_X1 g643(.A(new_n645_), .B1(new_n837_), .B2(KEYINPUT57), .C1(new_n843_), .C2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n837_), .A2(KEYINPUT57), .ZN(new_n846_));
  INV_X1    g645(.A(new_n842_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n823_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n848_), .B2(new_n646_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n836_), .A2(new_n845_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n296_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n813_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n594_), .A2(new_n623_), .A3(new_n663_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n319_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n813_), .B1(new_n850_), .B2(new_n657_), .ZN(new_n858_));
  OR3_X1    g657(.A1(new_n858_), .A2(KEYINPUT59), .A3(new_n854_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT59), .B1(new_n852_), .B2(new_n854_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n859_), .A2(new_n319_), .A3(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n857_), .B1(new_n861_), .B2(new_n856_), .ZN(G1340gat));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(KEYINPUT60), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n266_), .B2(KEYINPUT60), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n855_), .B(new_n867_), .C1(new_n866_), .C2(new_n865_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n859_), .A2(new_n265_), .A3(new_n860_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n863_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n855_), .A2(new_n871_), .A3(new_n697_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n859_), .A2(new_n296_), .A3(new_n860_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n871_), .ZN(G1342gat));
  INV_X1    g673(.A(G134gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n855_), .A2(new_n875_), .A3(new_n646_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n859_), .A2(new_n704_), .A3(new_n860_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n875_), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n663_), .A2(new_n593_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n725_), .A3(new_n623_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n852_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n319_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT120), .B(G141gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n265_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n697_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  OR2_X1    g688(.A1(new_n852_), .A2(new_n880_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G162gat), .B1(new_n890_), .B2(new_n703_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n852_), .A2(G162gat), .A3(new_n645_), .A4(new_n880_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(KEYINPUT121), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895_));
  INV_X1    g694(.A(G162gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n881_), .B2(new_n704_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n892_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n898_), .ZN(G1347gat));
  NOR3_X1   g698(.A1(new_n725_), .A2(new_n664_), .A3(new_n623_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n593_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n858_), .A2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(new_n504_), .A3(new_n319_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  INV_X1    g703(.A(G169gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n900_), .A2(new_n319_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT122), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n592_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n645_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n909_), .A2(new_n846_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n697_), .B1(new_n910_), .B2(new_n845_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n908_), .B1(new_n911_), .B2(new_n813_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n905_), .B1(new_n912_), .B2(KEYINPUT123), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n914_), .B(new_n908_), .C1(new_n911_), .C2(new_n813_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n904_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n908_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT123), .B1(new_n858_), .B2(new_n917_), .ZN(new_n918_));
  AND4_X1   g717(.A1(new_n904_), .A2(new_n918_), .A3(new_n915_), .A4(G169gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n903_), .B1(new_n916_), .B2(new_n919_), .ZN(G1348gat));
  NOR2_X1   g719(.A1(new_n852_), .A2(new_n901_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n266_), .A2(new_n505_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G176gat), .B1(new_n902_), .B2(new_n265_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n922_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(G1349gat));
  AOI21_X1  g726(.A(G183gat), .B1(new_n921_), .B2(new_n697_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n851_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n902_), .B2(new_n929_), .ZN(G1350gat));
  NAND4_X1  g729(.A1(new_n902_), .A2(new_n646_), .A3(new_n352_), .A4(new_n354_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n858_), .A2(new_n703_), .A3(new_n901_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n351_), .ZN(G1351gat));
  XNOR2_X1  g732(.A(KEYINPUT126), .B(G197gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n850_), .A2(new_n851_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n813_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n623_), .A2(new_n601_), .A3(new_n670_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n937_), .A2(KEYINPUT125), .A3(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n852_), .B2(new_n938_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n934_), .B1(new_n943_), .B2(new_n319_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n934_), .ZN(new_n945_));
  AOI211_X1 g744(.A(new_n661_), .B(new_n945_), .C1(new_n940_), .C2(new_n942_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1352gat));
  AOI21_X1  g746(.A(KEYINPUT125), .B1(new_n937_), .B2(new_n939_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n852_), .A2(new_n941_), .A3(new_n938_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n265_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(G204gat), .ZN(new_n951_));
  INV_X1    g750(.A(G204gat), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n943_), .A2(new_n952_), .A3(new_n265_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1353gat));
  OR2_X1    g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n943_), .B2(new_n296_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(KEYINPUT63), .B(G211gat), .ZN(new_n957_));
  AOI211_X1 g756(.A(new_n851_), .B(new_n957_), .C1(new_n940_), .C2(new_n942_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n958_), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n943_), .A2(new_n478_), .A3(new_n646_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n703_), .B1(new_n940_), .B2(new_n942_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n478_), .B2(new_n961_), .ZN(G1355gat));
endmodule


