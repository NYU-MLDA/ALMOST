//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n948_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_, new_n975_, new_n976_, new_n977_,
    new_n979_, new_n980_, new_n981_, new_n983_, new_n984_, new_n985_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n996_, new_n997_, new_n998_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT64), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n214_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n212_), .A2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n217_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT65), .A3(new_n217_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  AND3_X1   g031(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(new_n213_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n235_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT9), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n237_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n235_), .B1(new_n209_), .B2(new_n237_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n234_), .B(new_n236_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n222_), .B1(new_n232_), .B2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n210_), .B1(new_n221_), .B2(KEYINPUT67), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n234_), .A2(new_n244_), .A3(new_n220_), .A4(new_n218_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT8), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G57gat), .B(G64gat), .Z(new_n248_));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G57gat), .B(G64gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT68), .B(G71gat), .ZN(new_n253_));
  INV_X1    g052(.A(G78gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G71gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT68), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G71gat), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n257_), .A2(new_n259_), .A3(new_n254_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n250_), .B(new_n252_), .C1(new_n255_), .C2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n259_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G78gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n253_), .A2(new_n254_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT11), .A4(new_n251_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n205_), .B1(new_n247_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n221_), .A2(KEYINPUT67), .ZN(new_n268_));
  INV_X1    g067(.A(new_n210_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n245_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n211_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n214_), .A2(new_n219_), .A3(new_n236_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(new_n239_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n227_), .A2(new_n231_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n274_), .A2(new_n275_), .B1(new_n221_), .B2(new_n212_), .ZN(new_n276_));
  AOI211_X1 g075(.A(KEYINPUT12), .B(new_n266_), .C1(new_n271_), .C2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n276_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n261_), .A2(new_n265_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n267_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n242_), .B2(new_n246_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n271_), .A2(new_n276_), .A3(new_n266_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n205_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G120gat), .B(G148gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G204gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G176gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n282_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT69), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT69), .B1(new_n293_), .B2(new_n294_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n202_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n294_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT13), .A3(new_n295_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G29gat), .B(G50gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G43gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G36gat), .ZN(new_n308_));
  INV_X1    g107(.A(G36gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G43gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n306_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n309_), .A2(G43gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n307_), .A2(G36gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT71), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n305_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G15gat), .B(G22gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G1gat), .A2(G8gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT14), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G1gat), .ZN(new_n328_));
  INV_X1    g127(.A(G8gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n324_), .A2(new_n325_), .A3(new_n330_), .A4(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n314_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n323_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n323_), .A2(KEYINPUT79), .A3(new_n334_), .A4(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n332_), .A2(new_n333_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n320_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G229gat), .A2(G233gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n343_), .B(KEYINPUT80), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n340_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n334_), .A2(new_n319_), .A3(new_n314_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n342_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n343_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n342_), .A2(KEYINPUT78), .A3(new_n349_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G113gat), .B(G141gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G169gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G197gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n348_), .A2(new_n355_), .A3(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n346_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n358_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT81), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n341_), .B(KEYINPUT77), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G231gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(new_n280_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G127gat), .B(G155gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT16), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G183gat), .ZN(new_n376_));
  INV_X1    g175(.A(G211gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT17), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n373_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n379_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n373_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n304_), .A2(new_n369_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G127gat), .B(G134gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G113gat), .B(G120gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G183gat), .ZN(new_n393_));
  INV_X1    g192(.A(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n392_), .A2(new_n395_), .B1(G169gat), .B2(G176gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT22), .B(G169gat), .ZN(new_n397_));
  INV_X1    g196(.A(G176gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT83), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G169gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT22), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT22), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G169gat), .ZN(new_n403_));
  AND4_X1   g202(.A1(KEYINPUT83), .A2(new_n401_), .A3(new_n403_), .A4(new_n398_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n396_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT24), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n400_), .A3(new_n398_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G169gat), .A2(G176gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT24), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G169gat), .A2(G176gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n393_), .A2(KEYINPUT25), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT25), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G183gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n394_), .A2(KEYINPUT26), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT26), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G190gat), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT25), .B(G183gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G190gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(KEYINPUT82), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n417_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n405_), .A2(new_n430_), .A3(KEYINPUT30), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT30), .B1(new_n405_), .B2(new_n430_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G71gat), .B(G99gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n432_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n436_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n405_), .A2(new_n430_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n438_), .B1(new_n441_), .B2(new_n431_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n389_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n436_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n431_), .A3(new_n438_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n388_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G15gat), .B(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT31), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT29), .ZN(new_n454_));
  AND3_X1   g253(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT1), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT1), .ZN(new_n461_));
  NAND3_X1  g260(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G155gat), .A2(G162gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n457_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n469_));
  OAI22_X1  g268(.A1(new_n468_), .A2(new_n469_), .B1(G141gat), .B2(G148gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n465_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n469_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT2), .B1(new_n475_), .B2(new_n467_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n477_));
  INV_X1    g276(.A(G141gat), .ZN(new_n478_));
  INV_X1    g277(.A(G148gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n474_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n472_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n472_), .B2(new_n484_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n454_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G22gat), .B(G50gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT28), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n455_), .A2(new_n456_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n464_), .B1(new_n494_), .B2(new_n461_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n470_), .B1(new_n495_), .B2(new_n457_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n483_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT2), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n473_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT86), .B1(new_n496_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n486_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n454_), .A3(new_n491_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n493_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(KEYINPUT29), .A3(new_n486_), .ZN(new_n506_));
  INV_X1    g305(.A(G218gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G211gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n377_), .A2(G218gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT21), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G197gat), .B(G204gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT21), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n513_), .A2(KEYINPUT21), .A3(new_n508_), .A4(new_n509_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(G228gat), .A2(G233gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT29), .B1(new_n496_), .B2(new_n500_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n517_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n506_), .A2(new_n520_), .B1(new_n523_), .B2(new_n519_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n505_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n489_), .A2(new_n492_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n491_), .B1(new_n502_), .B2(new_n454_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT87), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G78gat), .B(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n493_), .A2(new_n503_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n529_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT87), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n525_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n531_), .B2(KEYINPUT87), .ZN(new_n535_));
  AOI211_X1 g334(.A(new_n504_), .B(new_n529_), .C1(new_n493_), .C2(new_n503_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n505_), .A2(new_n524_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n453_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n452_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n449_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n525_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n537_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n410_), .A2(new_n395_), .A3(new_n411_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n413_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n401_), .A2(new_n403_), .A3(KEYINPUT90), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT90), .B1(new_n401_), .B2(new_n403_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n548_), .B1(new_n551_), .B2(new_n398_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n424_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n553_), .A2(new_n416_), .A3(new_n412_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n522_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n405_), .A2(new_n430_), .A3(new_n517_), .A4(new_n516_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT20), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G226gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT19), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n558_), .B(KEYINPUT88), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT19), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n564_), .A3(KEYINPUT89), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n562_), .A2(new_n563_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n560_), .A2(KEYINPUT19), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n557_), .A2(new_n565_), .A3(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G64gat), .B(G92gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G8gat), .B(G36gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n402_), .A2(G169gat), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n400_), .A2(KEYINPUT22), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n401_), .A2(new_n403_), .A3(KEYINPUT90), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n398_), .A3(new_n582_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n396_), .A2(new_n583_), .B1(new_n417_), .B2(new_n424_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n577_), .B1(new_n584_), .B2(new_n518_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n439_), .A2(new_n522_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n567_), .A2(new_n568_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n570_), .A2(new_n576_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n569_), .A2(new_n565_), .ZN(new_n590_));
  AND4_X1   g389(.A1(KEYINPUT20), .A2(new_n555_), .A3(new_n590_), .A4(new_n556_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n587_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n575_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n593_), .A3(KEYINPUT27), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT94), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n589_), .A2(new_n593_), .A3(new_n596_), .A4(KEYINPUT27), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n599_));
  AND3_X1   g398(.A1(new_n570_), .A2(new_n576_), .A3(new_n588_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n576_), .B1(new_n570_), .B2(new_n588_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n472_), .A2(new_n484_), .A3(new_n388_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n472_), .A2(new_n484_), .A3(new_n388_), .A4(KEYINPUT92), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n501_), .A2(new_n389_), .A3(new_n486_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G225gat), .A2(G233gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G1gat), .B(G29gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT0), .ZN(new_n612_));
  INV_X1    g411(.A(G57gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(G85gat), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n607_), .A2(new_n608_), .A3(KEYINPUT4), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT4), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n501_), .A2(new_n617_), .A3(new_n389_), .A4(new_n486_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n609_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n610_), .B(new_n615_), .C1(new_n616_), .C2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n607_), .A2(new_n608_), .A3(KEYINPUT4), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n619_), .A3(new_n618_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n615_), .B1(new_n624_), .B2(new_n610_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n598_), .A2(new_n602_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT32), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n575_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT93), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(KEYINPUT93), .B(new_n630_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n570_), .B(new_n588_), .C1(new_n629_), .C2(new_n575_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n635_), .B(new_n636_), .C1(new_n622_), .C2(new_n625_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n621_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n600_), .A2(new_n601_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n624_), .A2(KEYINPUT33), .A3(new_n610_), .A4(new_n615_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n623_), .A2(new_n609_), .A3(new_n618_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n615_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n607_), .A2(new_n608_), .A3(new_n619_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .A4(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n637_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n453_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n648_));
  AOI22_X1  g447(.A1(new_n546_), .A2(new_n628_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(G190gat), .B(G218gat), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(G134gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT74), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(G162gat), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G162gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n652_), .B(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT36), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n279_), .A2(new_n335_), .A3(new_n323_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n247_), .A2(new_n320_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(G232gat), .A2(G233gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT34), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT35), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT70), .Z(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT73), .B1(new_n662_), .B2(KEYINPUT35), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n662_), .A2(KEYINPUT73), .A3(KEYINPUT35), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n664_), .A2(KEYINPUT75), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n659_), .A2(new_n660_), .A3(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n664_), .A2(KEYINPUT75), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n669_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n671_), .A2(new_n660_), .A3(new_n659_), .A4(new_n667_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n655_), .A2(new_n658_), .A3(new_n670_), .A4(new_n672_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n670_), .A2(new_n672_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n655_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n649_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n385_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n626_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G1gat), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT38), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT37), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n673_), .B2(KEYINPUT76), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n675_), .ZN(new_n685_));
  OAI221_X1 g484(.A(new_n673_), .B1(KEYINPUT76), .B2(new_n683_), .C1(new_n674_), .C2(new_n655_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n649_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n385_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT96), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n385_), .A2(new_n688_), .A3(KEYINPUT96), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n691_), .A2(new_n328_), .A3(new_n679_), .A4(new_n692_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(KEYINPUT97), .A3(new_n682_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT97), .B1(new_n693_), .B2(new_n682_), .ZN(new_n695_));
  OAI221_X1 g494(.A(new_n681_), .B1(new_n682_), .B2(new_n693_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT98), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1324gat));
  AND2_X1   g497(.A1(new_n598_), .A2(new_n602_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n329_), .B1(new_n678_), .B2(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT39), .Z(new_n702_));
  AND2_X1   g501(.A1(new_n691_), .A2(new_n692_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n699_), .A2(G8gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT99), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n703_), .A2(KEYINPUT99), .A3(new_n704_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT40), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(G1325gat));
  INV_X1    g508(.A(G15gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n703_), .A2(new_n710_), .A3(new_n453_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n711_), .A2(KEYINPUT100), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(KEYINPUT100), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n678_), .B2(new_n453_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT41), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n712_), .A2(new_n713_), .A3(new_n715_), .ZN(G1326gat));
  INV_X1    g515(.A(G22gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n534_), .A2(new_n538_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n678_), .B2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n703_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1327gat));
  NAND2_X1  g522(.A1(new_n647_), .A2(new_n648_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n543_), .A2(new_n544_), .B1(new_n452_), .B2(new_n451_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n727_), .B2(new_n627_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n676_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n303_), .A2(new_n368_), .A3(new_n384_), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n729_), .A2(KEYINPUT104), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n729_), .B2(new_n730_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G29gat), .B1(new_n733_), .B2(new_n679_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n627_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n647_), .A2(new_n648_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n735_), .B(new_n687_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT102), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n728_), .A2(new_n740_), .A3(new_n735_), .A4(new_n687_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n687_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n649_), .B2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n730_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(KEYINPUT44), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT103), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n744_), .A2(new_n748_), .A3(KEYINPUT44), .A4(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT44), .B1(new_n744_), .B2(new_n745_), .ZN(new_n751_));
  INV_X1    g550(.A(G29gat), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n626_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n734_), .B1(new_n750_), .B2(new_n753_), .ZN(G1328gat));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n751_), .A2(new_n699_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n309_), .B1(new_n750_), .B2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n731_), .A2(new_n309_), .A3(new_n700_), .A4(new_n732_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n755_), .B(KEYINPUT46), .C1(new_n757_), .C2(new_n760_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1329gat));
  NAND3_X1  g564(.A1(new_n731_), .A2(new_n453_), .A3(new_n732_), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT106), .B(G43gat), .Z(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n768_), .B(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n750_), .ZN(new_n771_));
  OR3_X1    g570(.A1(new_n751_), .A2(new_n307_), .A3(new_n542_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n770_), .B(new_n774_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1330gat));
  AOI21_X1  g577(.A(G50gat), .B1(new_n733_), .B2(new_n718_), .ZN(new_n779_));
  INV_X1    g578(.A(G50gat), .ZN(new_n780_));
  INV_X1    g579(.A(new_n718_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n751_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n779_), .B1(new_n750_), .B2(new_n782_), .ZN(G1331gat));
  NAND2_X1  g582(.A1(new_n304_), .A2(new_n369_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n784_), .A2(new_n384_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n688_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n613_), .A3(new_n679_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n677_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G57gat), .B1(new_n788_), .B2(new_n626_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1332gat));
  OAI21_X1  g589(.A(G64gat), .B1(new_n788_), .B2(new_n699_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT48), .ZN(new_n792_));
  INV_X1    g591(.A(G64gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n786_), .A2(new_n793_), .A3(new_n700_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1333gat));
  OAI21_X1  g594(.A(G71gat), .B1(new_n788_), .B2(new_n542_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT49), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n542_), .A2(G71gat), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT109), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n786_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(G1334gat));
  OAI21_X1  g600(.A(G78gat), .B1(new_n788_), .B2(new_n781_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n786_), .A2(new_n254_), .A3(new_n718_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1335gat));
  INV_X1    g605(.A(new_n384_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n784_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n744_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(G85gat), .B1(new_n809_), .B2(new_n626_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n676_), .A3(new_n728_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n206_), .A3(new_n679_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(G1336gat));
  OAI21_X1  g613(.A(G92gat), .B1(new_n809_), .B2(new_n699_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n207_), .A3(new_n700_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1337gat));
  NAND3_X1  g616(.A1(new_n744_), .A2(new_n453_), .A3(new_n808_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n453_), .A2(new_n230_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n818_), .A2(G99gat), .B1(new_n812_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(KEYINPUT113), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT113), .B1(new_n820_), .B2(new_n821_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n820_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT51), .B1(new_n820_), .B2(new_n824_), .ZN(new_n826_));
  OAI22_X1  g625(.A1(new_n822_), .A2(new_n823_), .B1(new_n825_), .B2(new_n826_), .ZN(G1338gat));
  NAND3_X1  g626(.A1(new_n812_), .A2(new_n217_), .A3(new_n718_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n744_), .A2(new_n718_), .A3(new_n808_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n217_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n828_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT53), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n828_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1339gat));
  NOR3_X1   g639(.A1(new_n700_), .A2(new_n539_), .A3(new_n626_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(KEYINPUT59), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n352_), .A2(new_n354_), .A3(new_n345_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n358_), .A3(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n846_), .A2(new_n360_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n301_), .A2(new_n295_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n284_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n205_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n282_), .A2(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n267_), .B(KEYINPUT55), .C1(new_n277_), .C2(new_n281_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n854_), .B2(new_n292_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n291_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n851_), .A2(new_n282_), .B1(new_n849_), .B2(new_n205_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n853_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n855_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n367_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n366_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n294_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n848_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n675_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n866_), .B2(KEYINPUT116), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n368_), .B(new_n294_), .C1(new_n855_), .C2(new_n860_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n676_), .B1(new_n870_), .B2(new_n848_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n868_), .B1(new_n869_), .B2(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n854_), .A2(new_n292_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n856_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n284_), .A2(new_n204_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n283_), .A2(KEYINPUT12), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n279_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n284_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n884_));
  OAI22_X1  g683(.A1(KEYINPUT55), .A2(new_n882_), .B1(new_n884_), .B2(new_n204_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n853_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n857_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT117), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n854_), .A2(new_n889_), .A3(new_n857_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n878_), .A2(new_n888_), .A3(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n847_), .A2(new_n294_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n876_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(KEYINPUT58), .A3(new_n892_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n687_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n807_), .B1(new_n874_), .B2(new_n896_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n687_), .A2(new_n384_), .A3(new_n368_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n303_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(new_n303_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n843_), .B1(new_n897_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n895_), .A2(new_n687_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n893_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n894_), .A2(KEYINPUT119), .A3(new_n687_), .A4(new_n895_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n871_), .A2(KEYINPUT57), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n867_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n910_));
  AOI211_X1 g709(.A(KEYINPUT116), .B(new_n676_), .C1(new_n870_), .C2(new_n848_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n384_), .B1(new_n908_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n902_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n842_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n903_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G113gat), .B1(new_n917_), .B2(new_n369_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n915_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n369_), .A2(G113gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1340gat));
  OAI211_X1 g720(.A(new_n903_), .B(new_n304_), .C1(new_n915_), .C2(new_n916_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(G120gat), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n303_), .A2(KEYINPUT60), .ZN(new_n924_));
  MUX2_X1   g723(.A(new_n924_), .B(KEYINPUT60), .S(G120gat), .Z(new_n925_));
  AND2_X1   g724(.A1(new_n906_), .A2(new_n907_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n807_), .B1(new_n926_), .B2(new_n874_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n841_), .B(new_n925_), .C1(new_n927_), .C2(new_n902_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n915_), .A2(KEYINPUT120), .A3(new_n925_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n923_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n923_), .A2(new_n932_), .A3(KEYINPUT121), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1341gat));
  OAI21_X1  g736(.A(G127gat), .B1(new_n917_), .B2(new_n384_), .ZN(new_n938_));
  OR2_X1    g737(.A1(new_n384_), .A2(G127gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n919_), .B2(new_n939_), .ZN(G1342gat));
  OAI21_X1  g739(.A(G134gat), .B1(new_n917_), .B2(new_n742_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n675_), .A2(G134gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n919_), .B2(new_n942_), .ZN(G1343gat));
  AOI21_X1  g742(.A(new_n545_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n944_), .A2(new_n679_), .A3(new_n699_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n369_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n478_), .ZN(G1344gat));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n303_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n479_), .ZN(G1345gat));
  NOR2_X1   g748(.A1(new_n945_), .A2(new_n384_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT61), .B(G155gat), .Z(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1346gat));
  OAI21_X1  g751(.A(G162gat), .B1(new_n945_), .B2(new_n742_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n676_), .A2(new_n656_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n945_), .B2(new_n954_), .ZN(G1347gat));
  XNOR2_X1  g754(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n699_), .A2(new_n679_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n726_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n368_), .B(new_n960_), .C1(new_n897_), .C2(new_n902_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n400_), .B1(new_n961_), .B2(KEYINPUT122), .ZN(new_n962_));
  INV_X1    g761(.A(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n961_), .A2(KEYINPUT122), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n957_), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n962_), .B(new_n956_), .C1(KEYINPUT122), .C2(new_n961_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n897_), .A2(new_n902_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n967_), .A2(new_n959_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n968_), .A2(new_n368_), .A3(new_n551_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n965_), .A2(new_n966_), .A3(new_n969_), .ZN(G1348gat));
  AOI21_X1  g769(.A(G176gat), .B1(new_n968_), .B2(new_n304_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n718_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n972_));
  AND4_X1   g771(.A1(G176gat), .A2(new_n304_), .A3(new_n453_), .A4(new_n958_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n971_), .B1(new_n972_), .B2(new_n973_), .ZN(G1349gat));
  INV_X1    g773(.A(new_n968_), .ZN(new_n975_));
  NOR3_X1   g774(.A1(new_n975_), .A2(new_n384_), .A3(new_n427_), .ZN(new_n976_));
  NAND4_X1  g775(.A1(new_n972_), .A2(new_n807_), .A3(new_n453_), .A4(new_n958_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n976_), .B1(new_n393_), .B2(new_n977_), .ZN(G1350gat));
  OAI21_X1  g777(.A(G190gat), .B1(new_n975_), .B2(new_n742_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n676_), .A2(new_n428_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(new_n980_), .B(KEYINPUT124), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n979_), .B1(new_n975_), .B2(new_n981_), .ZN(G1351gat));
  NAND2_X1  g781(.A1(new_n944_), .A2(new_n958_), .ZN(new_n983_));
  INV_X1    g782(.A(new_n983_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n984_), .A2(new_n368_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g785(.A1(new_n984_), .A2(new_n304_), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n987_), .B(G204gat), .ZN(G1353gat));
  OAI21_X1  g787(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n989_));
  AOI21_X1  g788(.A(new_n384_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n990_));
  INV_X1    g789(.A(new_n990_), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n989_), .B1(new_n983_), .B2(new_n991_), .ZN(new_n992_));
  NOR3_X1   g791(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n993_));
  XNOR2_X1  g792(.A(new_n993_), .B(KEYINPUT126), .ZN(new_n994_));
  XOR2_X1   g793(.A(new_n992_), .B(new_n994_), .Z(G1354gat));
  AOI21_X1  g794(.A(G218gat), .B1(new_n984_), .B2(new_n676_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n687_), .A2(G218gat), .ZN(new_n997_));
  XOR2_X1   g796(.A(new_n997_), .B(KEYINPUT127), .Z(new_n998_));
  AOI21_X1  g797(.A(new_n996_), .B1(new_n984_), .B2(new_n998_), .ZN(G1355gat));
endmodule


