//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203_));
  AND3_X1   g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT11), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n203_), .B1(new_n202_), .B2(KEYINPUT11), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  OAI22_X1  g009(.A1(new_n204_), .A2(new_n205_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(KEYINPUT65), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n221_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n228_));
  AND2_X1   g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n220_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n214_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT10), .B(G99gat), .Z(new_n237_));
  AOI22_X1  g036(.A1(new_n226_), .A2(new_n230_), .B1(new_n237_), .B2(new_n217_), .ZN(new_n238_));
  INV_X1    g037(.A(G85gat), .ZN(new_n239_));
  INV_X1    g038(.A(G92gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT9), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n241_), .A2(new_n242_), .B1(new_n243_), .B2(G92gat), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT9), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT64), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(new_n243_), .A3(new_n242_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n240_), .A2(KEYINPUT9), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n247_), .B(new_n248_), .C1(new_n234_), .C2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n238_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n218_), .A2(new_n219_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n229_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT8), .A3(new_n234_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n236_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n213_), .A2(KEYINPUT12), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n236_), .A2(new_n251_), .A3(new_n256_), .A4(KEYINPUT66), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n213_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT12), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n261_), .A2(new_n262_), .A3(new_n212_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(KEYINPUT68), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n261_), .A2(new_n272_), .A3(new_n262_), .A4(new_n212_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n264_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n268_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n274_), .A2(KEYINPUT69), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n274_), .B2(new_n275_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n270_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G120gat), .B(G148gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G176gat), .B(G204gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n270_), .B(new_n285_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n284_), .A2(KEYINPUT13), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT13), .B1(new_n284_), .B2(new_n286_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT71), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G29gat), .B(G36gat), .Z(new_n295_));
  XOR2_X1   g094(.A(G43gat), .B(G50gat), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G29gat), .B(G36gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G43gat), .B(G50gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n263_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n301_), .B(KEYINPUT15), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n257_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G232gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT34), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT35), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n303_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G190gat), .B(G218gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n305_), .A2(KEYINPUT72), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n257_), .A2(new_n304_), .A3(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n317_), .B(new_n319_), .C1(new_n263_), .C2(new_n302_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n308_), .A2(KEYINPUT35), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n320_), .A2(KEYINPUT73), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT73), .B1(new_n320_), .B2(new_n321_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n311_), .B(new_n316_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n321_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n320_), .A2(KEYINPUT73), .A3(new_n321_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n310_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n314_), .B(KEYINPUT36), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n324_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT75), .B1(new_n331_), .B2(KEYINPUT37), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(KEYINPUT75), .A3(KEYINPUT37), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT37), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n324_), .B(new_n335_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT76), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n311_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n330_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n335_), .A4(new_n324_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n333_), .A2(new_n334_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G8gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT77), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G15gat), .B(G22gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G1gat), .A2(G8gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT14), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n344_), .A2(KEYINPUT77), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n344_), .A2(KEYINPUT77), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n351_), .A2(new_n348_), .A3(new_n346_), .A4(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G231gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT78), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n354_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(new_n213_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G127gat), .B(G155gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT16), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G183gat), .B(G211gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT17), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n363_), .A2(new_n364_), .ZN(new_n366_));
  OR3_X1    g165(.A1(new_n359_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n359_), .A2(new_n365_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n343_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n294_), .A2(new_n371_), .A3(KEYINPUT79), .ZN(new_n372_));
  INV_X1    g171(.A(G197gat), .ZN(new_n373_));
  INV_X1    g172(.A(G204gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT87), .B(G197gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n374_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT21), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT89), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n373_), .A2(KEYINPUT87), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT87), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G197gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n383_), .A3(new_n374_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n378_), .B1(G197gat), .B2(G204gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n386_), .A2(KEYINPUT88), .ZN(new_n387_));
  XOR2_X1   g186(.A(G211gat), .B(G218gat), .Z(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n386_), .B2(KEYINPUT88), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n377_), .A2(new_n390_), .A3(new_n378_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n380_), .A2(new_n387_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n377_), .A2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(KEYINPUT90), .B(new_n375_), .C1(new_n376_), .C2(new_n374_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n395_), .A2(KEYINPUT21), .A3(new_n396_), .A4(new_n388_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n392_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT1), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT1), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G155gat), .A3(G162gat), .ZN(new_n404_));
  OR2_X1    g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .A4(KEYINPUT83), .ZN(new_n406_));
  XOR2_X1   g205(.A(G141gat), .B(G148gat), .Z(new_n407_));
  OAI211_X1 g206(.A(new_n406_), .B(new_n407_), .C1(KEYINPUT83), .C2(new_n404_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409_));
  INV_X1    g208(.A(G141gat), .ZN(new_n410_));
  INV_X1    g209(.A(G148gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n412_), .A2(new_n414_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n408_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n398_), .A2(new_n399_), .B1(new_n400_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(G228gat), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n408_), .A2(new_n418_), .A3(KEYINPUT84), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT84), .B1(new_n408_), .B2(new_n418_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(KEYINPUT85), .A3(KEYINPUT29), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n419_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n408_), .A2(new_n418_), .A3(KEYINPUT84), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT29), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n426_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n421_), .A2(new_n426_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G78gat), .B(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT92), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n400_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G22gat), .B(G50gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT28), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n443_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT85), .B1(new_n429_), .B2(KEYINPUT29), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n434_), .A2(new_n435_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n438_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n392_), .A2(new_n397_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT91), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n392_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n452_), .A2(new_n453_), .B1(KEYINPUT29), .B2(new_n419_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n450_), .B(new_n441_), .C1(new_n454_), .C2(new_n425_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n421_), .A2(new_n426_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n441_), .B1(new_n457_), .B2(new_n450_), .ZN(new_n458_));
  OAI22_X1  g257(.A1(new_n442_), .A2(new_n447_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n450_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n440_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n461_), .A2(KEYINPUT92), .A3(new_n455_), .A4(new_n446_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G183gat), .A2(G190gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT23), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(G183gat), .B2(G190gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G169gat), .A2(G176gat), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G176gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT22), .B(G169gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT93), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(new_n472_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n470_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(G169gat), .A2(G176gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(KEYINPUT24), .A3(new_n468_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n466_), .A2(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT25), .B(G183gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT26), .B(G190gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n476_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n451_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G226gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT19), .ZN(new_n488_));
  NOR2_X1   g287(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G169gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n467_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n392_), .A2(new_n397_), .A3(new_n484_), .A4(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n486_), .A2(KEYINPUT20), .A3(new_n488_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT20), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n484_), .A2(new_n491_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n451_), .B2(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n469_), .A2(new_n475_), .B1(new_n483_), .B2(new_n479_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n392_), .A3(new_n397_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n488_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G8gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G64gat), .B(G92gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n494_), .A2(new_n500_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n497_), .A2(new_n499_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n488_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n505_), .B1(new_n510_), .B2(new_n493_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n464_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n452_), .A2(new_n453_), .A3(new_n498_), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n451_), .B2(new_n496_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n509_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n486_), .A2(KEYINPUT20), .A3(new_n509_), .A4(new_n492_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n505_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n506_), .B1(new_n494_), .B2(new_n500_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(KEYINPUT27), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n512_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G127gat), .B(G134gat), .Z(new_n524_));
  XOR2_X1   g323(.A(G113gat), .B(G120gat), .Z(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT82), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G127gat), .B(G134gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G113gat), .B(G120gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n526_), .B1(new_n531_), .B2(KEYINPUT82), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n432_), .A2(new_n433_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G225gat), .A2(G233gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n420_), .A2(new_n531_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n432_), .A2(KEYINPUT95), .A3(new_n433_), .A4(new_n532_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT98), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n538_), .A2(new_n537_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n536_), .A4(new_n535_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G1gat), .B(G29gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT97), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G85gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n536_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT4), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n541_), .B2(new_n535_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n533_), .A2(new_n552_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n551_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n544_), .A2(new_n550_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n550_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n540_), .A2(new_n543_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT95), .B1(new_n429_), .B2(new_n532_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n538_), .A2(new_n537_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT4), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n536_), .B1(new_n562_), .B2(new_n554_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n559_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n532_), .B(KEYINPUT31), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G99gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G227gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(G15gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT30), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n572_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n484_), .B2(new_n491_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT81), .B(G43gat), .ZN(new_n575_));
  OR3_X1    g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n565_), .A2(new_n567_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n575_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n578_));
  AND4_X1   g377(.A1(new_n568_), .A2(new_n576_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n568_), .A2(new_n577_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n557_), .A2(new_n564_), .A3(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n463_), .A2(new_n523_), .A3(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n544_), .A2(new_n556_), .A3(KEYINPUT33), .A4(new_n550_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT99), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n559_), .A2(new_n563_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n587_), .A2(KEYINPUT99), .A3(KEYINPUT33), .A4(new_n550_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n557_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n510_), .A2(new_n493_), .A3(new_n505_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n521_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n551_), .B1(new_n562_), .B2(new_n554_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n541_), .A2(new_n551_), .A3(new_n535_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n558_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n586_), .A2(new_n588_), .A3(new_n590_), .A4(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n459_), .A2(new_n462_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n557_), .A2(new_n564_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n506_), .A2(KEYINPUT32), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n510_), .B2(new_n493_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n517_), .A2(new_n519_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n599_), .A3(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n512_), .A2(new_n522_), .A3(new_n564_), .A4(new_n557_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n581_), .B1(new_n607_), .B2(new_n463_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n583_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n354_), .A2(new_n301_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT80), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n354_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n302_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n612_), .B(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n304_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n616_), .A3(new_n610_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n618_), .A2(new_n620_), .A3(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n372_), .A2(new_n609_), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT79), .B1(new_n294_), .B2(new_n371_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AOI21_X1  g433(.A(G1gat), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n600_), .A2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n632_), .A2(KEYINPUT102), .A3(KEYINPUT38), .A4(new_n636_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n629_), .B(new_n369_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n638_));
  AND4_X1   g437(.A1(new_n588_), .A2(new_n586_), .A3(new_n590_), .A4(new_n597_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n605_), .A2(new_n462_), .A3(new_n459_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n608_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n583_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n331_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n331_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT103), .B1(new_n609_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n638_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n638_), .B2(new_n648_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n600_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G1gat), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n630_), .A2(new_n631_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n636_), .ZN(new_n655_));
  OAI22_X1  g454(.A1(new_n654_), .A2(new_n655_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n637_), .A2(new_n653_), .A3(new_n656_), .ZN(G1324gat));
  INV_X1    g456(.A(new_n523_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(G8gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n638_), .A2(new_n648_), .A3(new_n523_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G8gat), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(KEYINPUT39), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(KEYINPUT39), .ZN(new_n663_));
  OAI22_X1  g462(.A1(new_n654_), .A2(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(G1325gat));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n581_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(G15gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n668_), .B2(G15gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n672_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(KEYINPUT106), .A3(new_n670_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676_));
  INV_X1    g475(.A(new_n581_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(G15gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n632_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n678_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n654_), .A2(KEYINPUT107), .A3(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n673_), .B(new_n675_), .C1(new_n679_), .C2(new_n681_), .ZN(G1326gat));
  OR3_X1    g481(.A1(new_n654_), .A2(G22gat), .A3(new_n599_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n463_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(G22gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n684_), .B2(G22gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(G1327gat));
  NOR2_X1   g487(.A1(new_n609_), .A2(new_n629_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n646_), .A2(new_n369_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n293_), .A2(new_n689_), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n600_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n643_), .B(new_n343_), .C1(KEYINPUT108), .C2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n337_), .A2(new_n342_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n331_), .A2(KEYINPUT75), .A3(KEYINPUT37), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n697_), .B(KEYINPUT108), .C1(new_n332_), .C2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n332_), .B2(new_n698_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n699_), .B(KEYINPUT43), .C1(new_n609_), .C2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n696_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n369_), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n629_), .B(new_n703_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n702_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n702_), .B2(new_n704_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n600_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n694_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NOR3_X1   g508(.A1(new_n692_), .A2(G36gat), .A3(new_n658_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n705_), .A2(new_n706_), .A3(new_n658_), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(KEYINPUT110), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(KEYINPUT110), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n715_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  NAND2_X1  g520(.A1(new_n693_), .A2(new_n581_), .ZN(new_n722_));
  INV_X1    g521(.A(G43gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  NOR4_X1   g525(.A1(new_n705_), .A2(new_n706_), .A3(new_n723_), .A4(new_n677_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n726_), .A2(KEYINPUT47), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT47), .B1(new_n726_), .B2(new_n727_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1330gat));
  NOR2_X1   g529(.A1(new_n599_), .A2(G50gat), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT114), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n693_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n702_), .A2(new_n704_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n702_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .A4(new_n463_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(G50gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n736_), .A2(new_n463_), .A3(new_n738_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT112), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT113), .B1(new_n740_), .B2(new_n742_), .ZN(new_n743_));
  AND4_X1   g542(.A1(KEYINPUT113), .A2(new_n742_), .A3(G50gat), .A4(new_n739_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n733_), .B1(new_n743_), .B2(new_n744_), .ZN(G1331gat));
  NOR2_X1   g544(.A1(new_n369_), .A2(new_n628_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n648_), .A2(new_n294_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n600_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n294_), .A2(new_n643_), .A3(new_n629_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(new_n371_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n748_), .A2(G57gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1332gat));
  OAI21_X1  g553(.A(G64gat), .B1(new_n747_), .B2(new_n658_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT48), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n658_), .A2(G64gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n752_), .B2(new_n757_), .ZN(G1333gat));
  OR3_X1    g557(.A1(new_n752_), .A2(G71gat), .A3(new_n677_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n747_), .A2(new_n677_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G71gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G71gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1334gat));
  OAI21_X1  g563(.A(G78gat), .B1(new_n747_), .B2(new_n599_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT50), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n599_), .A2(G78gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n752_), .B2(new_n767_), .ZN(G1335gat));
  NOR2_X1   g567(.A1(new_n750_), .A2(new_n690_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n600_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT115), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n703_), .A2(new_n628_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n702_), .A2(new_n294_), .A3(new_n772_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n773_), .A2(new_n239_), .A3(new_n748_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n771_), .A2(new_n774_), .ZN(G1336gat));
  NAND3_X1  g574(.A1(new_n769_), .A2(new_n240_), .A3(new_n523_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G92gat), .B1(new_n773_), .B2(new_n658_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1337gat));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n581_), .A3(new_n237_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G99gat), .B1(new_n773_), .B2(new_n677_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n769_), .A2(new_n217_), .A3(new_n463_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  INV_X1    g583(.A(new_n773_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n463_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n786_), .B2(G106gat), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT52), .B(new_n217_), .C1(new_n785_), .C2(new_n463_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n783_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n783_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  AND2_X1   g592(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n616_), .B1(new_n354_), .B2(new_n301_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n624_), .B1(new_n619_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n615_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n617_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n627_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n212_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n258_), .B(new_n267_), .C1(new_n801_), .C2(KEYINPUT12), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n264_), .A2(new_n265_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n803_), .A2(new_n269_), .A3(new_n804_), .A4(new_n258_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n258_), .B1(new_n801_), .B2(KEYINPUT12), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n267_), .A2(new_n268_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT55), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AOI221_X4 g607(.A(KEYINPUT117), .B1(new_n275_), .B2(new_n802_), .C1(new_n805_), .C2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n805_), .A2(new_n808_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n802_), .A2(new_n275_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n283_), .B1(new_n809_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT56), .B(new_n283_), .C1(new_n809_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n286_), .A2(new_n628_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n286_), .A2(new_n628_), .A3(KEYINPUT116), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n800_), .B1(new_n818_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n794_), .B1(new_n824_), .B2(new_n646_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n794_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n821_), .A2(new_n822_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n817_), .B2(new_n816_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n331_), .B(new_n827_), .C1(new_n829_), .C2(new_n800_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n825_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n817_), .A2(KEYINPUT118), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n804_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n806_), .A2(KEYINPUT55), .A3(new_n807_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n812_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n811_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(KEYINPUT56), .A4(new_n283_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n832_), .A2(new_n840_), .A3(new_n816_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n286_), .A2(new_n627_), .A3(new_n798_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(KEYINPUT58), .A3(new_n842_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n343_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n703_), .B1(new_n831_), .B2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n700_), .A2(new_n289_), .A3(new_n746_), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT54), .Z(new_n850_));
  OR2_X1    g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n463_), .A2(new_n748_), .A3(new_n523_), .A4(new_n677_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n628_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(G113gat), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n852_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n852_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT59), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n858_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n628_), .A2(KEYINPUT121), .A3(G113gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(KEYINPUT121), .B2(G113gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n855_), .B1(new_n864_), .B2(new_n866_), .ZN(G1340gat));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n293_), .B2(KEYINPUT60), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n868_), .A2(KEYINPUT60), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n851_), .A2(new_n852_), .A3(new_n869_), .A4(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n857_), .A2(new_n294_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n868_), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n851_), .A2(new_n703_), .A3(new_n852_), .ZN(new_n875_));
  INV_X1    g674(.A(G127gat), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n369_), .A2(new_n876_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n864_), .B2(new_n878_), .ZN(G1342gat));
  NAND3_X1  g678(.A1(new_n851_), .A2(new_n646_), .A3(new_n852_), .ZN(new_n880_));
  INV_X1    g679(.A(G134gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n700_), .A2(new_n881_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n864_), .B2(new_n883_), .ZN(G1343gat));
  NOR2_X1   g683(.A1(new_n599_), .A2(new_n581_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n600_), .A3(new_n658_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT122), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n851_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n410_), .A3(new_n628_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G141gat), .B1(new_n888_), .B2(new_n629_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1344gat));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n411_), .A3(new_n294_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G148gat), .B1(new_n888_), .B2(new_n293_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1345gat));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  OR3_X1    g695(.A1(new_n888_), .A2(new_n369_), .A3(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n888_), .B2(new_n369_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n888_), .B2(new_n700_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n331_), .A2(G162gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n888_), .B2(new_n901_), .ZN(G1347gat));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n658_), .A2(new_n463_), .A3(new_n582_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n628_), .B(new_n904_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n905_), .B2(G169gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  INV_X1    g706(.A(new_n905_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n473_), .A2(new_n474_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n906_), .A2(new_n907_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n906_), .A2(new_n907_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n905_), .A2(new_n903_), .A3(G169gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1348gat));
  XNOR2_X1  g713(.A(KEYINPUT124), .B(G176gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n470_), .A2(KEYINPUT124), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n851_), .A2(new_n294_), .A3(new_n904_), .ZN(new_n917_));
  MUX2_X1   g716(.A(new_n915_), .B(new_n916_), .S(new_n917_), .Z(G1349gat));
  NAND2_X1  g717(.A1(new_n851_), .A2(new_n904_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920_));
  OAI22_X1  g719(.A1(new_n919_), .A2(new_n369_), .B1(new_n920_), .B2(G183gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n851_), .A2(new_n703_), .A3(new_n904_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n481_), .B1(KEYINPUT125), .B2(G183gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n919_), .B2(new_n700_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n646_), .A2(new_n482_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n919_), .B2(new_n926_), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n885_), .A2(new_n748_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n523_), .B1(new_n928_), .B2(KEYINPUT126), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(KEYINPUT126), .B2(new_n928_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n851_), .A2(new_n628_), .A3(new_n930_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g731(.A1(new_n851_), .A2(new_n294_), .A3(new_n930_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n851_), .A2(new_n703_), .A3(new_n930_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  OAI211_X1 g738(.A(new_n343_), .B(new_n930_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(G218gat), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n851_), .A2(new_n930_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n331_), .A2(G218gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n941_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(KEYINPUT127), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n946_), .B(new_n941_), .C1(new_n942_), .C2(new_n943_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1355gat));
endmodule


