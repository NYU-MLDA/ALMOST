//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G155gat), .ZN(new_n203_));
  INV_X1    g002(.A(G162gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT1), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G155gat), .A3(G162gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n205_), .B(new_n207_), .C1(G155gat), .C2(G162gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(G141gat), .B(G148gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT90), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT90), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n212_), .A3(new_n209_), .ZN(new_n213_));
  NOR3_X1   g012(.A1(KEYINPUT91), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n215_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G155gat), .B(G162gat), .Z(new_n221_));
  AOI22_X1  g020(.A1(new_n211_), .A2(new_n213_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT28), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G22gat), .B(G50gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT21), .ZN(new_n228_));
  AND2_X1   g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G197gat), .ZN(new_n232_));
  INV_X1    g031(.A(G204gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G197gat), .A2(G204gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(KEYINPUT21), .A3(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G218gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G211gat), .ZN(new_n240_));
  INV_X1    g039(.A(G211gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G218gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n243_), .A2(KEYINPUT21), .A3(new_n234_), .A4(new_n235_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n220_), .A2(new_n221_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n213_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n212_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n246_), .B1(new_n250_), .B2(KEYINPUT29), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT94), .ZN(new_n252_));
  INV_X1    g051(.A(G233gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n253_), .A2(KEYINPUT92), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(KEYINPUT92), .ZN(new_n255_));
  OAI21_X1  g054(.A(G228gat), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OR3_X1    g055(.A1(new_n251_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n252_), .B1(new_n251_), .B2(new_n256_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n238_), .A2(KEYINPUT93), .A3(new_n244_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT93), .B1(new_n238_), .B2(new_n244_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n256_), .B(new_n262_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT95), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n259_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n227_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n259_), .A2(new_n263_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n265_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n226_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n225_), .B(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n274_), .A3(new_n266_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G127gat), .B(G134gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT88), .ZN(new_n281_));
  XOR2_X1   g080(.A(G127gat), .B(G134gat), .Z(new_n282_));
  XOR2_X1   g081(.A(G113gat), .B(G120gat), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT89), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n250_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n280_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n247_), .B(new_n288_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G225gat), .A2(G233gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n281_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n289_), .B(KEYINPUT4), .C1(new_n293_), .C2(new_n222_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT100), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n287_), .A2(KEYINPUT100), .A3(KEYINPUT4), .A4(new_n289_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n290_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n287_), .B2(KEYINPUT4), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n292_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G1gat), .B(G29gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT101), .B(G85gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT0), .B(G57gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n300_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n307_), .B1(new_n310_), .B2(new_n292_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT22), .B(G169gat), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G183gat), .ZN(new_n318_));
  INV_X1    g117(.A(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT23), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n321_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(KEYINPUT83), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(G183gat), .A3(G190gat), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT23), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n320_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT97), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT97), .B(new_n320_), .C1(new_n326_), .C2(new_n330_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n317_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n337_));
  INV_X1    g136(.A(G169gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n314_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n339_), .A2(KEYINPUT24), .A3(new_n316_), .A4(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n318_), .A2(KEYINPUT25), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G183gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n319_), .A2(KEYINPUT26), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G190gat), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n342_), .A2(new_n344_), .A3(new_n345_), .A4(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n341_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT84), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(new_n321_), .B2(KEYINPUT23), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n352_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n327_), .A2(new_n329_), .A3(KEYINPUT23), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n338_), .A3(new_n314_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n349_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n336_), .A2(new_n246_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n339_), .A2(new_n340_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n357_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n341_), .A3(new_n348_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n326_), .A2(new_n330_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n354_), .A2(new_n355_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n367_), .A2(new_n368_), .B1(new_n369_), .B2(new_n317_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n364_), .B1(new_n262_), .B2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n360_), .A2(new_n363_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n359_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n245_), .B1(new_n335_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT98), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT98), .B(new_n245_), .C1(new_n335_), .C2(new_n373_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT96), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n327_), .A2(new_n329_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n324_), .B(new_n325_), .C1(new_n379_), .C2(KEYINPUT23), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n349_), .A3(new_n366_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n356_), .A2(new_n320_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n317_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n381_), .B(new_n384_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n378_), .B1(new_n385_), .B2(KEYINPUT20), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n378_), .B(KEYINPUT20), .C1(new_n262_), .C2(new_n370_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n376_), .B(new_n377_), .C1(new_n386_), .C2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n372_), .B1(new_n389_), .B2(new_n362_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT32), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT18), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n390_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT20), .B1(new_n262_), .B2(new_n370_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT96), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n387_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(new_n363_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n360_), .A2(new_n371_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n362_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(KEYINPUT32), .A3(new_n395_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n312_), .A2(new_n397_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT99), .B1(new_n390_), .B2(new_n395_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n376_), .A2(new_n377_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n388_), .A2(new_n386_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n362_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n372_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n396_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(KEYINPUT99), .A3(new_n396_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n302_), .B2(new_n308_), .ZN(new_n418_));
  NOR4_X1   g217(.A1(new_n310_), .A2(KEYINPUT33), .A3(new_n307_), .A4(new_n292_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n287_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n299_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n298_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n287_), .A2(new_n289_), .A3(new_n299_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n307_), .ZN(new_n425_));
  OAI22_X1  g224(.A1(new_n418_), .A2(new_n419_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n406_), .B1(new_n416_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT27), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n414_), .A2(new_n428_), .A3(new_n415_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n312_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n404_), .A2(new_n396_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT102), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n404_), .A2(KEYINPUT102), .A3(new_n396_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n428_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT103), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n434_), .A2(KEYINPUT103), .A3(new_n436_), .A4(new_n435_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n277_), .A2(new_n427_), .B1(new_n431_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G227gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT85), .ZN(new_n444_));
  INV_X1    g243(.A(G71gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G99gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G15gat), .B(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT86), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n447_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n370_), .B(KEYINPUT30), .Z(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT31), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n451_), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(new_n293_), .Z(new_n456_));
  OR2_X1    g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n456_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT104), .B1(new_n442_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n410_), .A2(new_n395_), .A3(new_n411_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT27), .ZN(new_n463_));
  AOI211_X1 g262(.A(new_n433_), .B(new_n395_), .C1(new_n401_), .C2(new_n403_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT103), .B1(new_n465_), .B2(new_n434_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n440_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n429_), .B(new_n430_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n426_), .B1(new_n415_), .B2(new_n414_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n406_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n277_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n460_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT104), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n459_), .A2(new_n312_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(new_n277_), .A3(new_n441_), .A4(new_n429_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n461_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT8), .ZN(new_n478_));
  XOR2_X1   g277(.A(G85gat), .B(G92gat), .Z(new_n479_));
  NOR2_X1   g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT66), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT66), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT65), .B1(new_n484_), .B2(new_n483_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n482_), .A2(new_n483_), .B1(new_n485_), .B2(new_n480_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT6), .Z(new_n488_));
  OAI21_X1  g287(.A(new_n479_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n489_), .B2(KEYINPUT67), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(KEYINPUT67), .B2(new_n489_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n488_), .B(KEYINPUT64), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n478_), .B(new_n479_), .C1(new_n492_), .C2(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n479_), .A2(KEYINPUT9), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n497_), .B(new_n498_), .C1(KEYINPUT9), .C2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n492_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n494_), .A2(KEYINPUT68), .A3(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT69), .B(G71gat), .ZN(new_n508_));
  INV_X1    g307(.A(G78gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n507_), .B1(new_n510_), .B2(KEYINPUT11), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n501_), .A2(KEYINPUT70), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n501_), .A2(KEYINPUT70), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n494_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT12), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n506_), .A2(new_n514_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n506_), .B2(new_n514_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G230gat), .A2(G233gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n522_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n506_), .A2(new_n514_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n513_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n520_), .A2(new_n521_), .A3(KEYINPUT71), .A4(new_n522_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n525_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G120gat), .B(G148gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G176gat), .B(G204gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n525_), .A2(new_n529_), .A3(new_n530_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT13), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(KEYINPUT13), .A3(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G29gat), .B(G36gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G15gat), .B(G22gat), .ZN(new_n550_));
  INV_X1    g349(.A(G8gat), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G1gat), .B(G8gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n547_), .B(KEYINPUT79), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n558_), .B(new_n556_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT80), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n564_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n544_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n477_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G127gat), .B(G155gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT76), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n556_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(new_n514_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n514_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT77), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n506_), .A2(new_n547_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT35), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT34), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n517_), .A2(new_n549_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT35), .A3(new_n590_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(KEYINPUT36), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n587_), .B(new_n592_), .C1(new_n588_), .C2(new_n591_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n594_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n599_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n597_), .B(KEYINPUT36), .Z(new_n602_));
  AND3_X1   g401(.A1(new_n601_), .A2(KEYINPUT75), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT75), .B1(new_n601_), .B2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n586_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n571_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT106), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n202_), .B1(new_n610_), .B2(new_n312_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n544_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n601_), .A2(new_n602_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n600_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT37), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT74), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n618_), .B(new_n600_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n612_), .A2(new_n585_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT78), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n569_), .ZN(new_n626_));
  AND4_X1   g425(.A1(new_n202_), .A2(new_n626_), .A3(new_n312_), .A4(new_n477_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT105), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n611_), .B1(new_n628_), .B2(KEYINPUT38), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(KEYINPUT38), .B2(new_n628_), .ZN(G1324gat));
  AND2_X1   g429(.A1(new_n626_), .A2(new_n477_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n441_), .A2(new_n429_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n551_), .A3(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n571_), .A2(new_n632_), .A3(new_n607_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(G8gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n634_), .B2(G8gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n633_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT108), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n633_), .B(new_n641_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n640_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1325gat));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n610_), .B2(new_n460_), .ZN(new_n648_));
  XOR2_X1   g447(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n649_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n631_), .A2(new_n647_), .A3(new_n460_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(G1326gat));
  OAI21_X1  g452(.A(G22gat), .B1(new_n609_), .B2(new_n277_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT42), .ZN(new_n655_));
  INV_X1    g454(.A(G22gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n631_), .A2(new_n656_), .A3(new_n276_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1327gat));
  NOR2_X1   g457(.A1(new_n585_), .A2(new_n605_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n571_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n661_), .B2(new_n312_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  INV_X1    g462(.A(new_n621_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n477_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT110), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n476_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT104), .B(new_n460_), .C1(new_n468_), .C2(new_n471_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n461_), .A2(KEYINPUT110), .A3(new_n474_), .A4(new_n476_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n664_), .A3(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT111), .B1(new_n671_), .B2(KEYINPUT43), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n665_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(KEYINPUT44), .A3(new_n586_), .A4(new_n570_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n675_), .A2(G29gat), .A3(new_n312_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n586_), .A3(new_n570_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n662_), .B1(new_n676_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  INV_X1    g480(.A(G36gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n632_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n570_), .A2(new_n586_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n671_), .A2(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n671_), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n684_), .B1(new_n689_), .B2(new_n665_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n683_), .B1(new_n690_), .B2(KEYINPUT44), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n682_), .B1(new_n691_), .B2(new_n679_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n661_), .A2(new_n682_), .A3(new_n632_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT45), .Z(new_n694_));
  OAI21_X1  g493(.A(new_n681_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n675_), .A2(new_n632_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n690_), .A2(KEYINPUT44), .ZN(new_n697_));
  OAI21_X1  g496(.A(G36gat), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n694_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(KEYINPUT46), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n695_), .A2(new_n700_), .ZN(G1329gat));
  AOI21_X1  g500(.A(G43gat), .B1(new_n661_), .B2(new_n460_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT112), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n675_), .A2(G43gat), .A3(new_n460_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n697_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT47), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n707_), .B(new_n703_), .C1(new_n704_), .C2(new_n697_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n661_), .B2(new_n276_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n675_), .A2(G50gat), .A3(new_n276_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n679_), .ZN(G1331gat));
  INV_X1    g511(.A(G57gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n612_), .A2(new_n568_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(new_n477_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n664_), .A2(new_n586_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n312_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n607_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n713_), .A3(new_n718_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n721_), .B2(KEYINPUT113), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(KEYINPUT113), .B2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g522(.A(G64gat), .B1(new_n720_), .B2(new_n683_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n683_), .A2(G64gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n717_), .B2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n720_), .B2(new_n459_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  INV_X1    g528(.A(new_n717_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n445_), .A3(new_n460_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1334gat));
  OAI21_X1  g531(.A(G78gat), .B1(new_n720_), .B2(new_n277_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(new_n509_), .A3(new_n276_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  INV_X1    g536(.A(G85gat), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n715_), .A2(new_n659_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n718_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT115), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n714_), .A2(new_n586_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n689_), .B2(new_n665_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n718_), .A2(new_n738_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(G1336gat));
  INV_X1    g544(.A(new_n739_), .ZN(new_n746_));
  INV_X1    g545(.A(G92gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n632_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n743_), .A2(new_n632_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n747_), .ZN(G1337gat));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(KEYINPUT51), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n460_), .A3(new_n495_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT116), .ZN(new_n754_));
  INV_X1    g553(.A(new_n742_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n674_), .A2(new_n460_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(G99gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n752_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n751_), .A2(KEYINPUT51), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n746_), .A2(new_n496_), .A3(new_n276_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n674_), .A2(new_n276_), .A3(new_n755_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G106gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G106gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT53), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n761_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1339gat));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n716_), .A2(new_n771_), .A3(new_n612_), .A4(new_n569_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT54), .B1(new_n622_), .B2(new_n568_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n563_), .A2(new_n567_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n562_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n560_), .B1(new_n558_), .B2(new_n555_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(new_n560_), .B1(new_n557_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n778_), .B2(new_n567_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n540_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT119), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n540_), .A2(new_n782_), .A3(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n539_), .A2(new_n568_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n525_), .A2(new_n786_), .A3(new_n530_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n520_), .A2(new_n521_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n526_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n523_), .A2(new_n786_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n526_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT118), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n787_), .A2(new_n790_), .A3(new_n791_), .A4(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n536_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n536_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n785_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n605_), .B1(new_n784_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n536_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n536_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n539_), .B(new_n779_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n621_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n797_), .A2(new_n798_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT58), .A3(new_n539_), .A4(new_n779_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n800_), .A2(new_n801_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n800_), .A2(new_n801_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n774_), .B1(new_n811_), .B2(new_n586_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n632_), .A2(new_n276_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n460_), .A3(new_n312_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n568_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n811_), .A2(new_n586_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n774_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n814_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(KEYINPUT59), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n569_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n817_), .B1(new_n825_), .B2(new_n816_), .ZN(G1340gat));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n827_));
  AOI21_X1  g626(.A(G120gat), .B1(new_n544_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n827_), .B2(G120gat), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n815_), .A2(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT120), .ZN(new_n831_));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n612_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(G1341gat));
  AOI21_X1  g633(.A(new_n585_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n585_), .B(new_n821_), .C1(new_n835_), .C2(new_n774_), .ZN(new_n836_));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(KEYINPUT121), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT121), .B1(new_n836_), .B2(new_n837_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n586_), .A2(new_n837_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT122), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT59), .B1(new_n820_), .B2(new_n821_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n812_), .A2(new_n823_), .A3(new_n814_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n841_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n847_), .B(new_n848_), .C1(new_n839_), .C2(new_n838_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n844_), .A2(new_n849_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n815_), .A2(new_n851_), .A3(new_n606_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n621_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(G1343gat));
  NOR3_X1   g653(.A1(new_n460_), .A2(new_n277_), .A3(new_n718_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n820_), .A2(new_n683_), .A3(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n569_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT123), .B(G141gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n856_), .A2(new_n612_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g660(.A1(new_n856_), .A2(new_n586_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  OAI21_X1  g663(.A(G162gat), .B1(new_n856_), .B2(new_n621_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n606_), .A2(new_n204_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n856_), .B2(new_n866_), .ZN(G1347gat));
  NOR2_X1   g666(.A1(new_n812_), .A2(new_n276_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n632_), .A2(new_n475_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n313_), .A3(new_n568_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n869_), .A2(new_n568_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT124), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n868_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n876_), .B2(G169gat), .ZN(new_n877_));
  AOI211_X1 g676(.A(KEYINPUT62), .B(new_n338_), .C1(new_n868_), .C2(new_n875_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n872_), .B1(new_n877_), .B2(new_n878_), .ZN(G1348gat));
  NOR2_X1   g678(.A1(new_n870_), .A2(new_n612_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n314_), .ZN(G1349gat));
  AOI21_X1  g680(.A(G183gat), .B1(new_n871_), .B2(new_n585_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n342_), .A2(new_n344_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n870_), .A2(new_n586_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1350gat));
  NAND4_X1  g684(.A1(new_n871_), .A2(new_n345_), .A3(new_n347_), .A4(new_n606_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n868_), .A2(new_n664_), .A3(new_n869_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT125), .B1(new_n887_), .B2(G190gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n886_), .B1(new_n889_), .B2(new_n890_), .ZN(G1351gat));
  AND3_X1   g690(.A1(new_n632_), .A2(new_n459_), .A3(new_n430_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n820_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n568_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n820_), .A2(new_n544_), .A3(new_n892_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(G204gat), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n820_), .A2(new_n899_), .A3(new_n544_), .A4(new_n892_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n233_), .B1(new_n897_), .B2(KEYINPUT126), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n903_));
  AND4_X1   g702(.A1(KEYINPUT127), .A2(new_n903_), .A3(G204gat), .A4(new_n900_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1353gat));
  NAND2_X1  g704(.A1(new_n893_), .A2(new_n585_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT63), .B(G211gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n906_), .B2(new_n909_), .ZN(G1354gat));
  NAND3_X1  g709(.A1(new_n893_), .A2(new_n239_), .A3(new_n606_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n893_), .A2(new_n664_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n239_), .ZN(G1355gat));
endmodule


