//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n969_, new_n970_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G92gat), .ZN(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT65), .ZN(new_n207_));
  OAI21_X1  g006(.A(G85gat), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT64), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n212_), .C1(G85gat), .C2(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(new_n206_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT10), .B(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(KEYINPUT6), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n220_), .A2(G106gat), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n218_), .A2(new_n219_), .A3(new_n226_), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n208_), .A2(new_n213_), .B1(KEYINPUT9), .B2(new_n216_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT66), .B1(new_n228_), .B2(new_n225_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  OR3_X1    g029(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n231_), .B(new_n232_), .C1(new_n222_), .C2(new_n224_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  XOR2_X1   g033(.A(G85gat), .B(G92gat), .Z(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n230_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n233_), .A2(new_n235_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT8), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n236_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n243_), .A2(new_n227_), .A3(new_n229_), .A4(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n240_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G57gat), .B(G64gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT11), .ZN(new_n249_));
  XOR2_X1   g048(.A(G71gat), .B(G78gat), .Z(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n248_), .A2(KEYINPUT11), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n203_), .B1(new_n247_), .B2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n240_), .A2(new_n245_), .A3(new_n255_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT69), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(KEYINPUT69), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n246_), .A2(KEYINPUT68), .A3(new_n254_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n242_), .A2(KEYINPUT70), .A3(new_n236_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n230_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n255_), .A2(KEYINPUT12), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n246_), .A2(new_n254_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n257_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n262_), .A3(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT5), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G176gat), .B(G204gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n264_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n264_), .B2(new_n276_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n202_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n284_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(KEYINPUT13), .A3(new_n282_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(KEYINPUT71), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(KEYINPUT71), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT74), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G43gat), .B(G50gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n293_), .A2(KEYINPUT74), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(KEYINPUT74), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n295_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302_));
  INV_X1    g101(.A(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(G8gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT14), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G8gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n297_), .A2(new_n300_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G229gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT80), .Z(new_n317_));
  INV_X1    g116(.A(KEYINPUT15), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n311_), .B(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n310_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(new_n309_), .A3(new_n314_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G113gat), .B(G141gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT81), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G169gat), .B(G197gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n317_), .A2(new_n321_), .A3(new_n326_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT83), .ZN(new_n331_));
  INV_X1    g130(.A(G169gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT22), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G176gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT22), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n342_));
  INV_X1    g141(.A(G183gat), .ZN(new_n343_));
  INV_X1    g142(.A(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n337_), .A2(new_n338_), .A3(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT25), .B(G183gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G190gat), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n348_), .A2(new_n349_), .A3(KEYINPUT82), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT82), .B1(new_n348_), .B2(new_n349_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT24), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n338_), .A2(KEYINPUT24), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n347_), .B1(new_n352_), .B2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G43gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n360_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G227gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(G15gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT30), .ZN(new_n369_));
  XOR2_X1   g168(.A(G127gat), .B(G134gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(G113gat), .B(G120gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n369_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n365_), .B(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(G155gat), .A3(G162gat), .ZN(new_n381_));
  INV_X1    g180(.A(G155gat), .ZN(new_n382_));
  INV_X1    g181(.A(G162gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n387_), .B2(KEYINPUT1), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n386_), .A3(KEYINPUT1), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n379_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n377_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n375_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n393_), .A2(new_n395_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n384_), .A2(new_n387_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n372_), .B1(new_n391_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n387_), .A2(KEYINPUT1), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT85), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n403_), .A2(new_n390_), .A3(new_n381_), .A4(new_n384_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n378_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G127gat), .B(G134gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(new_n371_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n398_), .A2(new_n399_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n401_), .A2(KEYINPUT4), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT96), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n401_), .A2(new_n409_), .A3(KEYINPUT96), .A4(KEYINPUT4), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n372_), .B(new_n415_), .C1(new_n391_), .C2(new_n400_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n401_), .A2(new_n409_), .A3(new_n417_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G85gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT0), .B(G57gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n422_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n419_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n422_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n426_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n374_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT103), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n356_), .A2(KEYINPUT92), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n357_), .B1(new_n356_), .B2(KEYINPUT92), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n355_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n344_), .A2(KEYINPUT26), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT26), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G190gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT91), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT91), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n349_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n446_), .A3(new_n348_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n439_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT93), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n338_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(KEYINPUT93), .A2(G169gat), .A3(G176gat), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n346_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n332_), .A2(KEYINPUT22), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n335_), .A2(G169gat), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT94), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT94), .B1(new_n453_), .B2(new_n454_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n334_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n448_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT21), .ZN(new_n460_));
  INV_X1    g259(.A(G197gat), .ZN(new_n461_));
  INV_X1    g260(.A(G204gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT87), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G204gat), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n461_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G197gat), .A2(G204gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n460_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G218gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(G211gat), .ZN(new_n470_));
  INV_X1    g269(.A(G211gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G218gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n463_), .A2(new_n465_), .A3(new_n461_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n460_), .B1(G197gat), .B2(G204gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n468_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n463_), .A2(new_n465_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n467_), .B1(new_n478_), .B2(G197gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n460_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n459_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n343_), .A2(KEYINPUT25), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G183gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n484_), .B1(new_n488_), .B2(new_n443_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n348_), .A2(new_n349_), .A3(KEYINPUT82), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n359_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n337_), .A2(new_n338_), .A3(new_n346_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n491_), .A2(new_n477_), .A3(new_n481_), .A4(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G226gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT19), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT90), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n483_), .A2(KEYINPUT20), .A3(new_n493_), .A4(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT98), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n491_), .A2(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n482_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n468_), .A2(new_n476_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n448_), .A3(new_n458_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(KEYINPUT20), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n495_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n360_), .B2(new_n502_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT98), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n483_), .A4(new_n497_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n499_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G8gat), .B(G36gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G64gat), .B(G92gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n493_), .A2(KEYINPUT20), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n502_), .B1(new_n448_), .B2(new_n458_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n496_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n495_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT20), .A4(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n522_), .A3(new_n515_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n523_), .A2(KEYINPUT27), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n517_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT100), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n497_), .B1(new_n507_), .B2(new_n483_), .ZN(new_n527_));
  AND4_X1   g326(.A1(KEYINPUT20), .A2(new_n501_), .A3(new_n521_), .A4(new_n503_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n516_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n523_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n526_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  AOI211_X1 g332(.A(KEYINPUT100), .B(new_n531_), .C1(new_n529_), .C2(new_n523_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n525_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT102), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n520_), .A2(new_n522_), .A3(new_n515_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n515_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n532_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT100), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n530_), .A2(new_n526_), .A3(new_n532_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT102), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n525_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G228gat), .A2(G233gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n549_), .B2(new_n502_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n404_), .A2(new_n378_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n482_), .B(new_n546_), .C1(new_n548_), .C2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G78gat), .B(G106gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT88), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n552_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n553_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G22gat), .B(G50gat), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n405_), .A2(new_n548_), .A3(new_n408_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n551_), .B2(new_n548_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n561_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n564_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n551_), .A2(new_n548_), .A3(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n560_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n550_), .A2(new_n552_), .A3(KEYINPUT89), .A4(new_n554_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n557_), .A2(new_n559_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n550_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n554_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n570_), .B(new_n567_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n436_), .B1(new_n545_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n577_), .ZN(new_n579_));
  AOI211_X1 g378(.A(KEYINPUT103), .B(new_n579_), .C1(new_n536_), .C2(new_n544_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n435_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n577_), .A2(new_n432_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n542_), .A2(new_n582_), .A3(new_n525_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n416_), .A2(new_n417_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n401_), .A2(new_n409_), .A3(new_n418_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n426_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n529_), .B(new_n523_), .C1(new_n585_), .C2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n430_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT33), .B1(new_n589_), .B2(new_n427_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(KEYINPUT33), .A3(new_n427_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n515_), .A2(KEYINPUT32), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n520_), .A2(new_n522_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT97), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n520_), .A2(new_n596_), .A3(new_n522_), .A4(new_n593_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n593_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n595_), .A2(new_n597_), .B1(new_n510_), .B2(new_n598_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n591_), .A2(new_n592_), .B1(new_n432_), .B2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n583_), .B1(new_n600_), .B2(new_n579_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n374_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT101), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n605_), .A3(new_n602_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n330_), .B1(new_n581_), .B2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n254_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(new_n611_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n310_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n610_), .A2(new_n611_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n308_), .A3(new_n612_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G183gat), .B(G211gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT17), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(KEYINPUT17), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n615_), .A2(new_n617_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT78), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n615_), .A2(new_n617_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n622_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT78), .B(new_n622_), .C1(new_n615_), .C2(new_n617_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT79), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n624_), .B(new_n632_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT35), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT75), .B1(new_n637_), .B2(new_n638_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n311_), .B(KEYINPUT15), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n230_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n311_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n644_), .A2(KEYINPUT73), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT73), .ZN(new_n647_));
  INV_X1    g446(.A(new_n641_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n319_), .B2(new_n270_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n246_), .A2(new_n301_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n640_), .B1(new_n646_), .B2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT73), .B1(new_n644_), .B2(new_n645_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(new_n650_), .A3(new_n647_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n639_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G134gat), .B(G162gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT36), .Z(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT76), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n652_), .A2(new_n655_), .A3(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n658_), .A2(KEYINPUT36), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT37), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n652_), .A2(new_n655_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n662_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n652_), .A2(new_n655_), .A3(new_n659_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT37), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n634_), .B1(new_n665_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n292_), .A2(new_n608_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n433_), .A2(G1gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT105), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n674_), .A2(new_n679_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT38), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n667_), .A2(new_n668_), .ZN(new_n684_));
  AOI221_X4 g483(.A(KEYINPUT102), .B1(new_n517_), .B2(new_n524_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n543_), .B1(new_n542_), .B2(new_n525_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n577_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT103), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n545_), .A2(new_n436_), .A3(new_n577_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n434_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n599_), .A2(new_n432_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n585_), .A2(new_n587_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT33), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n428_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n693_), .A2(new_n695_), .A3(new_n592_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n577_), .ZN(new_n698_));
  AOI211_X1 g497(.A(KEYINPUT101), .B(new_n374_), .C1(new_n698_), .C2(new_n583_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n605_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n684_), .B1(new_n690_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n634_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n288_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n330_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n581_), .A2(new_n607_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(KEYINPUT106), .A3(new_n684_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G1gat), .B1(new_n709_), .B2(new_n433_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n678_), .A2(KEYINPUT38), .A3(new_n680_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n683_), .A2(new_n710_), .A3(new_n711_), .ZN(G1324gat));
  INV_X1    g511(.A(new_n545_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n674_), .A2(new_n304_), .A3(new_n713_), .A4(new_n675_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n704_), .A2(new_n713_), .A3(new_n706_), .A4(new_n708_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(G8gat), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n715_), .B2(G8gat), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(KEYINPUT39), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT39), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n715_), .A2(G8gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT107), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n723_), .B2(new_n717_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n714_), .B1(new_n720_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT40), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT40), .B(new_n714_), .C1(new_n720_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1325gat));
  OAI21_X1  g528(.A(G15gat), .B1(new_n709_), .B2(new_n602_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT41), .Z(new_n731_));
  NAND2_X1  g530(.A1(new_n674_), .A2(new_n675_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n374_), .A2(new_n367_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(G1326gat));
  OAI21_X1  g533(.A(G22gat), .B1(new_n709_), .B2(new_n577_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT42), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n577_), .A2(G22gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n732_), .B2(new_n737_), .ZN(G1327gat));
  INV_X1    g537(.A(new_n684_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n634_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n705_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n608_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G29gat), .B1(new_n743_), .B2(new_n432_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n665_), .A2(new_n670_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n707_), .B2(new_n753_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n752_), .B(new_n749_), .C1(new_n581_), .C2(new_n607_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n706_), .A2(new_n634_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n747_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n707_), .A2(new_n753_), .A3(new_n748_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n752_), .B1(new_n581_), .B2(new_n607_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n751_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n757_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n745_), .A3(new_n746_), .A4(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n432_), .A2(G29gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n744_), .B1(new_n764_), .B2(new_n765_), .ZN(G1328gat));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n742_), .A2(G36gat), .A3(new_n545_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT45), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n756_), .A2(new_n747_), .A3(new_n757_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n761_), .A2(new_n762_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n713_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n769_), .B1(new_n772_), .B2(G36gat), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n767_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(G36gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n764_), .B2(new_n713_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT110), .B(KEYINPUT46), .C1(new_n777_), .C2(new_n769_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n775_), .A2(new_n778_), .ZN(G1329gat));
  NOR3_X1   g578(.A1(new_n742_), .A2(G43gat), .A3(new_n602_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n764_), .A2(new_n374_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(G43gat), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g582(.A(G50gat), .B1(new_n743_), .B2(new_n579_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n579_), .A2(G50gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n764_), .B2(new_n785_), .ZN(G1331gat));
  NAND2_X1  g585(.A1(new_n328_), .A2(new_n329_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n581_), .B2(new_n607_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n788_), .A2(new_n705_), .A3(new_n671_), .ZN(new_n789_));
  INV_X1    g588(.A(G57gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n432_), .ZN(new_n791_));
  AND4_X1   g590(.A1(new_n330_), .A2(new_n704_), .A3(new_n291_), .A4(new_n708_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(new_n432_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n793_), .B2(new_n790_), .ZN(G1332gat));
  INV_X1    g593(.A(G64gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n789_), .A2(new_n795_), .A3(new_n713_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n792_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G64gat), .B1(new_n797_), .B2(new_n545_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(KEYINPUT48), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(KEYINPUT48), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(G1333gat));
  INV_X1    g600(.A(G71gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n789_), .A2(new_n802_), .A3(new_n374_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G71gat), .B1(new_n797_), .B2(new_n602_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(KEYINPUT49), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(KEYINPUT49), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n803_), .B1(new_n805_), .B2(new_n806_), .ZN(G1334gat));
  INV_X1    g606(.A(G78gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n789_), .A2(new_n808_), .A3(new_n579_), .ZN(new_n809_));
  OAI21_X1  g608(.A(G78gat), .B1(new_n797_), .B2(new_n577_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(KEYINPUT50), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(KEYINPUT50), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n811_), .B2(new_n812_), .ZN(G1335gat));
  AOI21_X1  g612(.A(new_n740_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n788_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(new_n215_), .A3(new_n432_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n634_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n288_), .A2(new_n787_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n761_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT111), .B1(new_n761_), .B2(new_n819_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n822_), .A2(new_n433_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n817_), .B1(new_n824_), .B2(new_n215_), .ZN(G1336gat));
  OAI21_X1  g624(.A(new_n713_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT112), .Z(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n822_), .A2(new_n823_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G92gat), .B1(new_n816_), .B2(new_n713_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT113), .ZN(G1337gat));
  NOR3_X1   g631(.A1(new_n815_), .A2(new_n602_), .A3(new_n220_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n834_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n835_), .A2(new_n836_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n837_));
  OR2_X1    g636(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n838_));
  OAI21_X1  g637(.A(G99gat), .B1(new_n820_), .B2(new_n602_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1338gat));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n579_), .B(new_n819_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n844_), .A2(new_n845_), .A3(G106gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n844_), .B2(G106gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n843_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n844_), .A2(G106gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT116), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n844_), .A2(new_n845_), .A3(G106gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(KEYINPUT52), .A3(new_n851_), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n815_), .A2(G106gat), .A3(new_n577_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1339gat));
  AOI21_X1  g655(.A(new_n262_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n276_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n273_), .A2(KEYINPUT55), .A3(new_n262_), .A4(new_n275_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n280_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT56), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n281_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n863_), .A2(new_n787_), .A3(new_n282_), .A4(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n320_), .A2(new_n309_), .A3(new_n315_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n326_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n329_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n739_), .B1(new_n867_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT57), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n282_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n877_));
  AOI211_X1 g676(.A(KEYINPUT56), .B(new_n281_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n877_), .A2(new_n330_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n873_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n684_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(KEYINPUT118), .A3(new_n882_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n863_), .A2(new_n282_), .A3(new_n872_), .A4(new_n866_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT119), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n752_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n877_), .A2(new_n871_), .A3(new_n878_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(KEYINPUT58), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n886_), .A2(new_n887_), .A3(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n876_), .A2(new_n883_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n634_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n818_), .A2(new_n752_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n285_), .A2(new_n287_), .A3(new_n330_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT54), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n671_), .A2(new_n288_), .A3(new_n897_), .A4(new_n330_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n896_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n893_), .A2(new_n900_), .ZN(new_n901_));
  AOI211_X1 g700(.A(new_n433_), .B(new_n602_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(G113gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n787_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n907_), .A2(KEYINPUT120), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(KEYINPUT120), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n904_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n903_), .A2(KEYINPUT120), .A3(new_n907_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n330_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n906_), .B1(new_n912_), .B2(new_n905_), .ZN(G1340gat));
  INV_X1    g712(.A(G120gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n288_), .B2(KEYINPUT60), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n904_), .B(new_n915_), .C1(KEYINPUT60), .C2(new_n914_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n292_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n914_), .ZN(G1341gat));
  INV_X1    g717(.A(G127gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n904_), .A2(new_n919_), .A3(new_n818_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n634_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n919_), .ZN(G1342gat));
  INV_X1    g721(.A(G134gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n904_), .A2(new_n923_), .A3(new_n739_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n752_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(G1343gat));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n713_), .A2(new_n577_), .A3(new_n433_), .A4(new_n374_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n901_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n899_), .B1(new_n892_), .B2(new_n634_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n928_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT121), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n787_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT122), .B(G141gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1344gat));
  NAND2_X1  g735(.A1(new_n933_), .A2(new_n291_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(new_n933_), .B2(new_n818_), .ZN(new_n940_));
  AOI211_X1 g739(.A(KEYINPUT123), .B(new_n634_), .C1(new_n929_), .C2(new_n932_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT61), .B(G155gat), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n940_), .A2(new_n941_), .A3(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n927_), .B1(new_n901_), .B2(new_n928_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n930_), .A2(KEYINPUT121), .A3(new_n931_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n818_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(KEYINPUT123), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n933_), .A2(new_n939_), .A3(new_n818_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n942_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n944_), .A2(new_n950_), .ZN(G1346gat));
  INV_X1    g750(.A(new_n933_), .ZN(new_n952_));
  OAI21_X1  g751(.A(G162gat), .B1(new_n952_), .B2(new_n752_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n933_), .A2(new_n383_), .A3(new_n739_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1347gat));
  NAND2_X1  g754(.A1(new_n713_), .A2(new_n435_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(KEYINPUT124), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n930_), .A2(new_n579_), .A3(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n787_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n455_), .A2(new_n456_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n959_), .A2(G169gat), .ZN(new_n962_));
  XNOR2_X1  g761(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n961_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n964_), .B1(new_n962_), .B2(new_n963_), .ZN(G1348gat));
  NAND3_X1  g764(.A1(new_n958_), .A2(new_n334_), .A3(new_n705_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n958_), .A2(new_n291_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n967_), .B2(new_n334_), .ZN(G1349gat));
  NAND2_X1  g767(.A1(new_n958_), .A2(new_n818_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n969_), .A2(new_n348_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n970_), .B1(new_n343_), .B2(new_n969_), .ZN(G1350gat));
  NAND4_X1  g770(.A1(new_n958_), .A2(new_n444_), .A3(new_n446_), .A4(new_n739_), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n958_), .A2(new_n753_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n973_), .B2(new_n344_), .ZN(G1351gat));
  NOR4_X1   g773(.A1(new_n545_), .A2(new_n577_), .A3(new_n432_), .A4(new_n374_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n901_), .A2(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n901_), .A2(KEYINPUT126), .A3(new_n975_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n980_), .A2(new_n787_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g781(.A(new_n478_), .ZN(new_n983_));
  AND3_X1   g782(.A1(new_n901_), .A2(KEYINPUT126), .A3(new_n975_), .ZN(new_n984_));
  AOI21_X1  g783(.A(KEYINPUT126), .B1(new_n901_), .B2(new_n975_), .ZN(new_n985_));
  OAI211_X1 g784(.A(new_n983_), .B(new_n291_), .C1(new_n984_), .C2(new_n985_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(new_n986_), .A2(KEYINPUT127), .ZN(new_n987_));
  AND2_X1   g786(.A1(new_n986_), .A2(KEYINPUT127), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n980_), .A2(new_n291_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n989_), .A2(G204gat), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n987_), .B1(new_n988_), .B2(new_n990_), .ZN(G1353gat));
  AOI21_X1  g790(.A(new_n634_), .B1(new_n978_), .B2(new_n979_), .ZN(new_n992_));
  OR2_X1    g791(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n993_));
  NOR2_X1   g792(.A1(new_n992_), .A2(new_n993_), .ZN(new_n994_));
  XOR2_X1   g793(.A(KEYINPUT63), .B(G211gat), .Z(new_n995_));
  AOI21_X1  g794(.A(new_n994_), .B1(new_n992_), .B2(new_n995_), .ZN(G1354gat));
  NAND3_X1  g795(.A1(new_n980_), .A2(new_n469_), .A3(new_n739_), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n752_), .B1(new_n978_), .B2(new_n979_), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n997_), .B1(new_n998_), .B2(new_n469_), .ZN(G1355gat));
endmodule


