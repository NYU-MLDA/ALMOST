//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_;
  OR2_X1    g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n203_));
  AND2_X1   g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n205_));
  NAND4_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT89), .A4(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT89), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(new_n204_), .B2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n202_), .B(new_n206_), .C1(new_n210_), .C2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT90), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT87), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT22), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G169gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n219_), .A2(new_n221_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT88), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT87), .B(G176gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT88), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n217_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT89), .B1(new_n209_), .B2(KEYINPUT23), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT85), .B(KEYINPUT23), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(new_n209_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n202_), .A4(new_n206_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n215_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n209_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT86), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n234_), .B2(new_n209_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n243_), .B2(new_n240_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT84), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(G169gat), .B2(G176gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT24), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n248_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n247_), .A2(G169gat), .A3(G176gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n217_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n249_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G183gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT83), .B1(new_n256_), .B2(KEYINPUT25), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(G190gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n257_), .B(new_n258_), .C1(new_n259_), .C2(KEYINPUT83), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n244_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n238_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G71gat), .B(G99gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G43gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n262_), .B(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G127gat), .B(G134gat), .Z(new_n266_));
  XOR2_X1   g065(.A(G113gat), .B(G120gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270_));
  INV_X1    g069(.A(G15gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT30), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT31), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(new_n268_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n269_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n268_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281_));
  INV_X1    g080(.A(G141gat), .ZN(new_n282_));
  INV_X1    g081(.A(G148gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n290_), .A2(KEYINPUT92), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT92), .B1(new_n290_), .B2(new_n294_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n285_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n291_), .B1(new_n293_), .B2(KEYINPUT1), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n302_), .A2(KEYINPUT91), .B1(new_n303_), .B2(new_n292_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT91), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n305_), .B(new_n291_), .C1(new_n293_), .C2(KEYINPUT1), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n301_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n280_), .B1(new_n297_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n290_), .A2(new_n294_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT92), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n290_), .A2(KEYINPUT92), .A3(new_n294_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n302_), .A2(KEYINPUT91), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n292_), .A2(new_n303_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n306_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n300_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n268_), .A3(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n308_), .A2(KEYINPUT4), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT4), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n320_), .B(new_n280_), .C1(new_n297_), .C2(new_n307_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT98), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n317_), .B1(new_n296_), .B2(new_n295_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n324_), .A2(KEYINPUT98), .A3(new_n320_), .A4(new_n280_), .ZN(new_n325_));
  AND4_X1   g124(.A1(new_n279_), .A2(new_n319_), .A3(new_n323_), .A4(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n279_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n308_), .A2(new_n327_), .A3(new_n318_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G85gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT0), .B(G57gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT33), .B1(new_n326_), .B2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n319_), .A2(new_n323_), .A3(new_n327_), .A4(new_n325_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n308_), .A2(new_n279_), .A3(new_n318_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT99), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT99), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n308_), .A2(new_n318_), .A3(new_n339_), .A4(new_n279_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n335_), .A2(new_n336_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n226_), .A2(new_n216_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n244_), .B2(new_n202_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT96), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n206_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(new_n249_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n249_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(KEYINPUT96), .A3(new_n235_), .A4(new_n206_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n252_), .A2(new_n254_), .B1(new_n259_), .B2(new_n258_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n345_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G211gat), .B(G218gat), .Z(new_n354_));
  INV_X1    g153(.A(G204gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT94), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT94), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G204gat), .ZN(new_n358_));
  INV_X1    g157(.A(G197gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT21), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(G197gat), .B2(G204gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n354_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n359_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n361_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n364_), .A2(new_n365_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G211gat), .B(G218gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(new_n361_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n363_), .A2(new_n366_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n343_), .B1(new_n353_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT97), .ZN(new_n375_));
  INV_X1    g174(.A(new_n370_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n262_), .B2(new_n376_), .ZN(new_n377_));
  AOI211_X1 g176(.A(KEYINPUT97), .B(new_n370_), .C1(new_n238_), .C2(new_n261_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n371_), .B(new_n374_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n353_), .A2(new_n370_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT20), .B1(new_n262_), .B2(new_n376_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n373_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT18), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n379_), .A2(new_n387_), .A3(new_n382_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n338_), .A2(new_n340_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n392_), .A2(KEYINPUT33), .A3(new_n336_), .A4(new_n335_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n342_), .A2(new_n389_), .A3(new_n390_), .A4(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(KEYINPUT32), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n380_), .A2(new_n381_), .A3(new_n373_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n377_), .A2(new_n378_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n353_), .A2(new_n370_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT20), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n373_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n400_), .B2(KEYINPUT100), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT100), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n402_), .B(new_n373_), .C1(new_n397_), .C2(new_n399_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n395_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n335_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n332_), .B1(new_n405_), .B2(new_n391_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n341_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n379_), .A2(new_n395_), .A3(new_n382_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n394_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT95), .B(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n324_), .B2(KEYINPUT29), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415_));
  INV_X1    g214(.A(new_n413_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n313_), .A2(new_n415_), .A3(new_n317_), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n415_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G22gat), .B(G50gat), .Z(new_n420_));
  NOR3_X1   g219(.A1(new_n419_), .A2(new_n370_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n420_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT29), .B1(new_n297_), .B2(new_n307_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n376_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n418_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n420_), .B1(new_n419_), .B2(new_n370_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n376_), .A3(new_n422_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n417_), .A4(new_n414_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G228gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(G78gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n425_), .A2(new_n428_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n412_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n418_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n426_), .A2(new_n427_), .B1(new_n417_), .B2(new_n414_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n425_), .A2(new_n428_), .A3(new_n432_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n411_), .A3(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n410_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n407_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n389_), .A2(new_n390_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n387_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n390_), .A2(KEYINPUT27), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n443_), .B(new_n446_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n278_), .B1(new_n442_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n407_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n441_), .A2(new_n451_), .A3(new_n278_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n400_), .A2(KEYINPUT100), .ZN(new_n453_));
  INV_X1    g252(.A(new_n396_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n403_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n448_), .B1(new_n455_), .B2(new_n388_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT27), .B1(new_n389_), .B2(new_n390_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT101), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT101), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n446_), .B(new_n459_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n452_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n450_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(KEYINPUT9), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470_));
  OR2_X1    g269(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n471_));
  INV_X1    g270(.A(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  INV_X1    g274(.A(G92gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(KEYINPUT9), .A3(new_n463_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n469_), .A2(new_n470_), .A3(new_n474_), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n466_), .A2(new_n468_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n463_), .A2(KEYINPUT9), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT64), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n472_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT65), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n490_), .A2(new_n485_), .A3(new_n486_), .A4(new_n472_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n488_), .A2(new_n481_), .A3(new_n489_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n477_), .A2(new_n463_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n479_), .B(new_n484_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G29gat), .B(G36gat), .Z(new_n498_));
  XOR2_X1   g297(.A(G43gat), .B(G50gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G232gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT34), .ZN(new_n503_));
  OAI22_X1  g302(.A1(new_n497_), .A2(new_n501_), .B1(KEYINPUT35), .B2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n500_), .B(KEYINPUT15), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n492_), .A2(new_n494_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT8), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n484_), .A2(new_n510_), .A3(new_n479_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n484_), .B2(new_n479_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n504_), .B1(new_n505_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n503_), .A2(KEYINPUT35), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT76), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n514_), .B(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G190gat), .B(G218gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT77), .ZN(new_n519_));
  XOR2_X1   g318(.A(G134gat), .B(G162gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT36), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n521_), .B(KEYINPUT36), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n517_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n462_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT105), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n484_), .A2(new_n479_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT68), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n484_), .A2(new_n510_), .A3(new_n479_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n534_), .A2(new_n535_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n538_));
  XOR2_X1   g337(.A(G71gat), .B(G78gat), .Z(new_n539_));
  OR2_X1    g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n539_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT12), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT69), .B1(new_n536_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(new_n497_), .B2(new_n544_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n497_), .A2(new_n544_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n513_), .A2(new_n551_), .A3(KEYINPUT12), .A4(new_n544_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n546_), .A2(new_n550_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT67), .ZN(new_n555_));
  INV_X1    g354(.A(new_n553_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n533_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n509_), .A2(new_n557_), .A3(KEYINPUT66), .A4(new_n543_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n549_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n533_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT66), .B1(new_n560_), .B2(new_n543_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n555_), .B(new_n556_), .C1(new_n559_), .C2(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n554_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n556_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT67), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G120gat), .B(G148gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT72), .ZN(new_n568_));
  XOR2_X1   g367(.A(G176gat), .B(G204gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT73), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n566_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n575_));
  NAND4_X1  g374(.A1(new_n565_), .A2(new_n572_), .A3(new_n554_), .A4(new_n562_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n576_), .A2(KEYINPUT74), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(KEYINPUT74), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n574_), .B(new_n575_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n563_), .A2(new_n580_), .A3(new_n572_), .A4(new_n565_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(KEYINPUT74), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n581_), .A2(new_n582_), .B1(new_n566_), .B2(new_n573_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT13), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n579_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G15gat), .B(G22gat), .ZN(new_n587_));
  INV_X1    g386(.A(G1gat), .ZN(new_n588_));
  INV_X1    g387(.A(G8gat), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT14), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G1gat), .B(G8gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n592_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n591_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(KEYINPUT82), .A3(new_n500_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT82), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n595_), .A2(new_n599_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n501_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n601_), .A2(new_n604_), .B1(new_n501_), .B2(new_n603_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n601_), .A2(new_n604_), .B1(new_n505_), .B2(new_n603_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n608_), .B(new_n615_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n586_), .A2(KEYINPUT104), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT104), .B1(new_n586_), .B2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n543_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(new_n603_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G127gat), .B(G155gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT17), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n622_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n627_), .B(KEYINPUT17), .Z(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n622_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n618_), .A2(new_n619_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n532_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT106), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT106), .B1(new_n532_), .B2(new_n633_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G1gat), .B1(new_n638_), .B2(new_n451_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n586_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n528_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(new_n524_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n641_), .B2(new_n524_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n632_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n462_), .B2(new_n617_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n462_), .A2(new_n648_), .A3(new_n617_), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n640_), .B(new_n647_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n407_), .B(KEYINPUT103), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n588_), .A3(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT38), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n639_), .A2(new_n655_), .ZN(G1324gat));
  NAND2_X1  g455(.A1(new_n458_), .A2(new_n460_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n589_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G8gat), .B1(new_n634_), .B2(new_n657_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(KEYINPUT39), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(KEYINPUT39), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT40), .B(new_n659_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  NAND3_X1  g466(.A1(new_n652_), .A2(new_n271_), .A3(new_n278_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n278_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n669_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(new_n669_), .B2(G15gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n441_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n652_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(G22gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n676_), .B2(G22gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(G1327gat));
  NOR2_X1   g479(.A1(new_n530_), .A2(new_n631_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n586_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G29gat), .B1(new_n683_), .B2(new_n407_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n618_), .A2(new_n619_), .A3(new_n631_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n645_), .B1(new_n450_), .B2(new_n461_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n688_), .B(new_n645_), .C1(new_n450_), .C2(new_n461_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n685_), .A2(KEYINPUT107), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n579_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n581_), .A2(new_n582_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n585_), .B1(new_n692_), .B2(new_n574_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n617_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n586_), .A2(KEYINPUT104), .A3(new_n617_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n632_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT44), .B1(new_n690_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(G29gat), .A3(new_n653_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n687_), .A2(new_n689_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n696_), .A2(KEYINPUT107), .A3(new_n632_), .A4(new_n697_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n700_), .A2(new_n704_), .A3(KEYINPUT44), .A4(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n690_), .A2(new_n708_), .A3(KEYINPUT44), .A4(new_n700_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n684_), .B1(new_n703_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n657_), .A2(G36gat), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n683_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT109), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n683_), .A2(new_n716_), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(KEYINPUT45), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(G36gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n701_), .B1(new_n707_), .B2(new_n709_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n658_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n712_), .B1(new_n722_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n725_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n727_), .A2(KEYINPUT46), .A3(new_n721_), .A4(new_n720_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1329gat));
  INV_X1    g528(.A(G43gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n683_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n278_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n730_), .ZN(new_n734_));
  AND4_X1   g533(.A1(KEYINPUT110), .A2(new_n710_), .A3(new_n702_), .A4(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT110), .B1(new_n724_), .B2(new_n734_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n733_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT47), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n739_), .B(new_n733_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1330gat));
  INV_X1    g540(.A(new_n724_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G50gat), .B1(new_n742_), .B2(new_n441_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n441_), .A2(G50gat), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT111), .Z(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n731_), .B2(new_n745_), .ZN(G1331gat));
  NOR3_X1   g545(.A1(new_n586_), .A2(new_n632_), .A3(new_n617_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n532_), .A2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n451_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n617_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n462_), .A2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n647_), .A2(new_n586_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n653_), .ZN(new_n754_));
  OR3_X1    g553(.A1(new_n753_), .A2(G57gat), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n749_), .A2(new_n755_), .ZN(G1332gat));
  OAI21_X1  g555(.A(G64gat), .B1(new_n748_), .B2(new_n657_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n657_), .A2(G64gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n753_), .B2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n748_), .B2(new_n732_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n732_), .A2(G71gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n753_), .B2(new_n764_), .ZN(G1334gat));
  NAND4_X1  g564(.A1(new_n751_), .A2(new_n752_), .A3(new_n430_), .A4(new_n674_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G78gat), .B1(new_n748_), .B2(new_n441_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT50), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(KEYINPUT50), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT113), .B(new_n766_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1335gat));
  AND4_X1   g573(.A1(new_n632_), .A2(new_n704_), .A3(new_n750_), .A4(new_n640_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(new_n407_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n751_), .A2(new_n640_), .A3(new_n681_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n653_), .A2(new_n475_), .ZN(new_n778_));
  OAI22_X1  g577(.A1(new_n776_), .A2(new_n475_), .B1(new_n777_), .B2(new_n778_), .ZN(G1336gat));
  NOR3_X1   g578(.A1(new_n777_), .A2(G92gat), .A3(new_n657_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n775_), .A2(new_n658_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(G92gat), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT114), .ZN(G1337gat));
  NAND3_X1  g582(.A1(new_n278_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n777_), .A2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT116), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n775_), .A2(new_n278_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(G99gat), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT115), .B(new_n486_), .C1(new_n775_), .C2(new_n278_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR3_X1   g591(.A1(new_n777_), .A2(G106gat), .A3(new_n441_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n775_), .A2(new_n674_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n472_), .B1(new_n796_), .B2(KEYINPUT52), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n796_), .A2(KEYINPUT52), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n795_), .B(new_n797_), .C1(new_n796_), .C2(KEYINPUT52), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g602(.A1(new_n692_), .A2(new_n617_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n554_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n546_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n807_), .A2(KEYINPUT119), .A3(new_n556_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT119), .B1(new_n807_), .B2(new_n556_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n806_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n546_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(KEYINPUT55), .A4(new_n553_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT120), .B1(new_n554_), .B2(new_n805_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n573_), .B1(new_n810_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT56), .B(new_n573_), .C1(new_n810_), .C2(new_n815_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n804_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n609_), .A2(new_n607_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n615_), .C1(new_n607_), .C2(new_n605_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n614_), .A2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n583_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n530_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT57), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n692_), .A2(new_n614_), .A3(new_n822_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n645_), .B1(new_n828_), .B2(KEYINPUT58), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(KEYINPUT58), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT121), .B(new_n645_), .C1(new_n828_), .C2(KEYINPUT58), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n631_), .B1(new_n826_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n646_), .A2(new_n750_), .A3(new_n586_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT54), .Z(new_n837_));
  NOR2_X1   g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n674_), .A2(new_n732_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n658_), .A2(new_n840_), .A3(new_n754_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n838_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n617_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n836_), .B(KEYINPUT54), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n826_), .A2(new_n834_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n631_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT59), .A3(new_n841_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n838_), .B2(new_n842_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n750_), .A2(KEYINPUT122), .ZN(new_n852_));
  MUX2_X1   g651(.A(KEYINPUT122), .B(new_n852_), .S(G113gat), .Z(new_n853_));
  AOI21_X1  g652(.A(new_n844_), .B1(new_n851_), .B2(new_n853_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n586_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n843_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n586_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n855_), .ZN(G1341gat));
  XOR2_X1   g658(.A(KEYINPUT124), .B(G127gat), .Z(new_n860_));
  NOR2_X1   g659(.A1(new_n632_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n851_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n631_), .B(new_n841_), .C1(new_n835_), .C2(new_n837_), .ZN(new_n864_));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT123), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n864_), .A2(KEYINPUT123), .A3(new_n865_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n862_), .B(new_n863_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n866_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n861_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT125), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n872_), .ZN(G1342gat));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n843_), .A2(new_n874_), .A3(new_n529_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n645_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n874_), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n838_), .A2(new_n278_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(new_n674_), .A3(new_n657_), .A4(new_n653_), .ZN(new_n880_));
  OR3_X1    g679(.A1(new_n880_), .A2(G141gat), .A3(new_n750_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G141gat), .B1(new_n880_), .B2(new_n750_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1344gat));
  OR3_X1    g682(.A1(new_n880_), .A2(G148gat), .A3(new_n586_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G148gat), .B1(new_n880_), .B2(new_n586_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1345gat));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  OR3_X1    g686(.A1(new_n880_), .A2(new_n632_), .A3(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n880_), .B2(new_n632_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n880_), .B2(new_n876_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n530_), .A2(G162gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n880_), .B2(new_n892_), .ZN(G1347gat));
  NOR3_X1   g692(.A1(new_n840_), .A2(new_n657_), .A3(new_n653_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n847_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n222_), .B1(new_n895_), .B2(new_n617_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n895_), .A2(new_n229_), .A3(new_n617_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n900_), .B(new_n901_), .C1(new_n896_), .C2(new_n898_), .ZN(G1348gat));
  NAND2_X1  g701(.A1(new_n895_), .A2(new_n640_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n218_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n228_), .B2(new_n903_), .ZN(G1349gat));
  NAND2_X1  g704(.A1(new_n847_), .A2(new_n894_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n632_), .ZN(new_n907_));
  MUX2_X1   g706(.A(G183gat), .B(new_n259_), .S(new_n907_), .Z(G1350gat));
  NAND3_X1  g707(.A1(new_n895_), .A2(new_n258_), .A3(new_n529_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G190gat), .B1(new_n906_), .B2(new_n876_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1351gat));
  NOR3_X1   g710(.A1(new_n657_), .A2(new_n407_), .A3(new_n441_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n879_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n750_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT127), .B(G197gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1352gat));
  INV_X1    g715(.A(new_n913_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G204gat), .B1(new_n917_), .B2(new_n640_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n356_), .A2(new_n358_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n913_), .A2(new_n586_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1353gat));
  XOR2_X1   g720(.A(KEYINPUT63), .B(G211gat), .Z(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n631_), .A3(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n913_), .B2(new_n632_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1354gat));
  OAI21_X1  g725(.A(G218gat), .B1(new_n913_), .B2(new_n876_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n530_), .A2(G218gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n913_), .B2(new_n928_), .ZN(G1355gat));
endmodule


