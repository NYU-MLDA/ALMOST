//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n980_, new_n981_, new_n983_, new_n984_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n996_, new_n997_, new_n998_;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G211gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT16), .B(G183gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(G15gat), .A2(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G15gat), .A2(G22gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(G8gat), .A3(new_n211_), .ZN(new_n212_));
  AOI221_X4 g011(.A(G8gat), .B1(new_n206_), .B2(new_n207_), .C1(new_n212_), .C2(KEYINPUT14), .ZN(new_n213_));
  INV_X1    g012(.A(G8gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(KEYINPUT14), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n206_), .A2(new_n207_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT75), .B(G1gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n213_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221_));
  AND2_X1   g020(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n221_), .B1(new_n224_), .B2(G8gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n216_), .ZN(new_n226_));
  OAI21_X1  g025(.A(G8gat), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n215_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n218_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n220_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G231gat), .A2(G233gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n219_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n227_), .A2(new_n218_), .A3(new_n228_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G231gat), .A3(G233gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G71gat), .B(G78gat), .ZN(new_n241_));
  OR3_X1    g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n241_), .A3(KEYINPUT11), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT76), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n237_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n237_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n205_), .B1(new_n248_), .B2(KEYINPUT17), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(KEYINPUT77), .A3(new_n247_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n205_), .A2(KEYINPUT17), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G190gat), .B(G218gat), .Z(new_n256_));
  XOR2_X1   g055(.A(G134gat), .B(G162gat), .Z(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT36), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT72), .Z(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT73), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT73), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G99gat), .A2(G106gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT7), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT6), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(G99gat), .A3(G106gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT8), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G85gat), .B(G92gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n272_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n268_), .A2(new_n270_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n274_), .B1(new_n280_), .B2(new_n266_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n276_), .B1(new_n281_), .B2(new_n273_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT70), .B(G29gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G43gat), .ZN(new_n285_));
  INV_X1    g084(.A(G50gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G36gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G43gat), .A2(G50gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n288_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n284_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n292_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(new_n283_), .A3(new_n290_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G106gat), .ZN(new_n298_));
  INV_X1    g097(.A(G99gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT10), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT10), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G99gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n298_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT66), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n301_), .A2(G99gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n299_), .A2(KEYINPUT10), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT65), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n298_), .ZN(new_n314_));
  INV_X1    g113(.A(G85gat), .ZN(new_n315_));
  INV_X1    g114(.A(G92gat), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n315_), .A2(new_n316_), .A3(KEYINPUT9), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n275_), .A2(KEYINPUT9), .B1(new_n268_), .B2(new_n270_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n307_), .A2(new_n314_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n282_), .A2(new_n297_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n271_), .A2(KEYINPUT67), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n268_), .A2(new_n270_), .A3(new_n277_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n266_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n273_), .B1(new_n325_), .B2(new_n275_), .ZN(new_n326_));
  AOI211_X1 g125(.A(KEYINPUT8), .B(new_n274_), .C1(new_n266_), .C2(new_n271_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT68), .B1(new_n322_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n282_), .A2(new_n330_), .A3(new_n320_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n296_), .B(KEYINPUT15), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT71), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n336_));
  AOI211_X1 g135(.A(new_n336_), .B(new_n333_), .C1(new_n329_), .C2(new_n331_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n321_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G232gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT34), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(KEYINPUT35), .A3(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n282_), .A2(new_n330_), .A3(new_n320_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n330_), .B1(new_n282_), .B2(new_n320_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n334_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n336_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n332_), .A2(KEYINPUT71), .A3(new_n334_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n340_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT35), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n349_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n347_), .A2(new_n351_), .A3(new_n352_), .A4(new_n321_), .ZN(new_n353_));
  AOI211_X1 g152(.A(new_n261_), .B(new_n264_), .C1(new_n341_), .C2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n258_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(KEYINPUT36), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n341_), .A2(new_n356_), .A3(new_n353_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT37), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n262_), .B1(new_n341_), .B2(new_n353_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT37), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n341_), .A2(new_n356_), .A3(new_n353_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n255_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(G155gat), .B2(G162gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n367_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(G155gat), .A3(G162gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n370_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT1), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n375_), .A3(KEYINPUT90), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT89), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT89), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(G141gat), .A3(G148gat), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT2), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n386_), .B(new_n389_), .C1(KEYINPUT3), .C2(new_n378_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT91), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n384_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G113gat), .B(G120gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT87), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT4), .B1(new_n396_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n384_), .A2(new_n394_), .A3(new_n391_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n394_), .B1(new_n384_), .B2(new_n391_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n400_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n392_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(KEYINPUT98), .A3(new_n399_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT98), .ZN(new_n410_));
  INV_X1    g209(.A(new_n399_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n392_), .B2(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n402_), .B(new_n404_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n403_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G1gat), .B(G29gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(new_n315_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT0), .B(G57gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  AND3_X1   g220(.A1(new_n415_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n244_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT12), .B(new_n426_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G230gat), .A2(G233gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT64), .Z(new_n429_));
  OAI21_X1  g228(.A(new_n320_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT12), .B1(new_n430_), .B2(new_n426_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n426_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n427_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n429_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n432_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n430_), .A2(new_n426_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G120gat), .B(G148gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G204gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT5), .B(G176gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n434_), .A2(new_n438_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n444_), .B(new_n446_), .C1(KEYINPUT69), .C2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n334_), .A2(new_n230_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G229gat), .A2(G233gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT79), .B1(new_n235_), .B2(new_n297_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT79), .ZN(new_n457_));
  AOI211_X1 g256(.A(new_n457_), .B(new_n296_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n454_), .B(new_n455_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n230_), .A2(new_n296_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n455_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G141gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G169gat), .B(G197gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n459_), .A2(new_n463_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n453_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT27), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT19), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G204gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT93), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G204gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(G197gat), .ZN(new_n483_));
  INV_X1    g282(.A(G197gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(G204gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G211gat), .B(G218gat), .Z(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(KEYINPUT21), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT21), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT93), .B(G204gat), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n490_), .B(new_n485_), .C1(new_n491_), .C2(new_n484_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n483_), .A2(KEYINPUT94), .A3(new_n490_), .A4(new_n485_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G197gat), .A2(G204gat), .ZN(new_n497_));
  OAI211_X1 g296(.A(KEYINPUT21), .B(new_n497_), .C1(new_n491_), .C2(G197gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n487_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT95), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n487_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(KEYINPUT95), .A3(new_n498_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n489_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT25), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n506_), .A2(KEYINPUT80), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(KEYINPUT80), .ZN(new_n508_));
  OAI21_X1  g307(.A(G183gat), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT81), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT26), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G190gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT83), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT82), .B(G190gat), .ZN(new_n516_));
  INV_X1    g315(.A(G183gat), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n516_), .A2(KEYINPUT26), .B1(KEYINPUT25), .B2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT81), .B(G183gat), .C1(new_n507_), .C2(new_n508_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n511_), .A2(new_n515_), .A3(new_n518_), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G183gat), .A2(G190gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT23), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT23), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(G183gat), .A3(G190gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G169gat), .A2(G176gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT24), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n525_), .A2(KEYINPUT84), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT84), .B1(new_n525_), .B2(new_n528_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(G169gat), .A2(G176gat), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n532_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n520_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT85), .B(G176gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT22), .B(G169gat), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n532_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n516_), .A2(new_n517_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n525_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT20), .B1(new_n505_), .B2(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n503_), .A2(KEYINPUT95), .A3(new_n498_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT95), .B1(new_n503_), .B2(new_n498_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n488_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n525_), .A2(new_n528_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT96), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT25), .B(G183gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT26), .B(G190gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(KEYINPUT96), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n548_), .A2(new_n551_), .A3(new_n552_), .A4(new_n533_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n525_), .B1(G183gat), .B2(G190gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n537_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n546_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n477_), .B1(new_n543_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT20), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n546_), .B2(new_n556_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n505_), .A2(new_n542_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n476_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G64gat), .B(G92gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G8gat), .B(G36gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n558_), .A2(new_n562_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n474_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n558_), .A2(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n567_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n560_), .A2(new_n477_), .A3(new_n561_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n559_), .B1(new_n546_), .B2(new_n541_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n556_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n505_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n477_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n568_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n579_), .A3(KEYINPUT27), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n571_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G78gat), .B(G106gat), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT29), .B1(new_n405_), .B2(new_n406_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G228gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT92), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n546_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n408_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n584_), .B1(new_n546_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n582_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n405_), .A2(new_n406_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT28), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n593_), .A3(new_n587_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n393_), .A2(new_n587_), .A3(new_n395_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT28), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G22gat), .B(G50gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n593_), .B1(new_n592_), .B2(new_n587_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n595_), .A2(KEYINPUT28), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n584_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n505_), .B2(new_n588_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n546_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n582_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n591_), .A2(new_n599_), .A3(new_n602_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n602_), .A2(new_n599_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n604_), .A2(new_n606_), .A3(new_n605_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n606_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G15gat), .B(G43gat), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT30), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n534_), .A2(new_n615_), .A3(new_n540_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n534_), .B2(new_n540_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n614_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n541_), .A2(KEYINPUT30), .ZN(new_n619_));
  INV_X1    g418(.A(new_n614_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n534_), .A2(new_n615_), .A3(new_n540_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G227gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT86), .ZN(new_n624_));
  INV_X1    g423(.A(G71gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(G99gat), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n618_), .A2(new_n622_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT88), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n627_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n616_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n620_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT88), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n618_), .A2(new_n622_), .A3(new_n627_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n400_), .B(KEYINPUT31), .Z(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n630_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT88), .B(new_n638_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n613_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n581_), .A2(new_n643_), .A3(KEYINPUT101), .A4(new_n424_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n571_), .A2(new_n580_), .A3(new_n424_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n608_), .A2(new_n612_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n641_), .A3(new_n640_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n645_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n644_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n642_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n646_), .B2(new_n613_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n567_), .A2(KEYINPUT32), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n572_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n574_), .A2(new_n578_), .ZN(new_n655_));
  OAI221_X1 g454(.A(new_n654_), .B1(new_n655_), .B2(new_n653_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT99), .B1(new_n423_), .B2(KEYINPUT33), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n659_));
  INV_X1    g458(.A(new_n417_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n401_), .B1(new_n416_), .B2(KEYINPUT4), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n404_), .B2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n658_), .B(new_n659_), .C1(new_n662_), .C2(new_n421_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n657_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n415_), .A2(new_n417_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n421_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(KEYINPUT33), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n402_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(KEYINPUT100), .A3(new_n403_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n661_), .B2(new_n404_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n666_), .B1(new_n413_), .B2(new_n404_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n558_), .A2(new_n562_), .A3(new_n568_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n667_), .A2(new_n673_), .A3(new_n573_), .A4(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n656_), .B(new_n647_), .C1(new_n664_), .C2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n652_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n650_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n366_), .A2(new_n425_), .A3(new_n473_), .A4(new_n678_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n679_), .A2(KEYINPUT102), .A3(new_n224_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT102), .B1(new_n679_), .B2(new_n224_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT38), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n649_), .A2(new_n644_), .B1(new_n652_), .B2(new_n676_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n357_), .A2(new_n359_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n687_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n678_), .A2(KEYINPUT103), .A3(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n688_), .A2(new_n690_), .A3(new_n473_), .A4(new_n254_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G1gat), .B1(new_n691_), .B2(new_n424_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n680_), .A2(KEYINPUT38), .A3(new_n681_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT104), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n684_), .A2(new_n696_), .A3(new_n692_), .A4(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1324gat));
  AND2_X1   g497(.A1(new_n366_), .A2(new_n678_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n581_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(new_n214_), .A3(new_n473_), .A4(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G8gat), .B1(new_n691_), .B2(new_n581_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT105), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT39), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n705_), .B(G8gat), .C1(new_n691_), .C2(new_n581_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n703_), .A2(new_n704_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n701_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT40), .B(new_n701_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1325gat));
  OR2_X1    g512(.A1(new_n691_), .A2(new_n642_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT41), .B1(new_n714_), .B2(G15gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n699_), .A2(new_n473_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n642_), .A2(G15gat), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n716_), .A2(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(G1326gat));
  OR3_X1    g519(.A1(new_n718_), .A2(G22gat), .A3(new_n647_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G22gat), .B1(new_n691_), .B2(new_n647_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT106), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(G22gat), .C1(new_n691_), .C2(new_n647_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n723_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n724_), .B1(new_n723_), .B2(new_n726_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n721_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(KEYINPUT107), .B(new_n721_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1327gat));
  NOR3_X1   g532(.A1(new_n453_), .A2(new_n472_), .A3(new_n254_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n358_), .A2(new_n363_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n678_), .B2(new_n737_), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT43), .B(new_n736_), .C1(new_n650_), .C2(new_n677_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n734_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(KEYINPUT44), .B(new_n734_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G29gat), .B1(new_n744_), .B2(new_n424_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n678_), .A2(new_n687_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n734_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n424_), .A2(G29gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT108), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n745_), .A2(new_n751_), .ZN(G1328gat));
  NAND3_X1  g551(.A1(new_n742_), .A2(new_n700_), .A3(new_n743_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT109), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n742_), .A2(new_n755_), .A3(new_n700_), .A4(new_n743_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(G36gat), .A3(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n748_), .A2(new_n288_), .A3(new_n700_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT45), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n757_), .A2(KEYINPUT46), .A3(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1329gat));
  NAND3_X1  g563(.A1(new_n748_), .A2(new_n285_), .A3(new_n651_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n744_), .A2(new_n642_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n285_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(G1330gat));
  OAI21_X1  g568(.A(G50gat), .B1(new_n744_), .B2(new_n647_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n748_), .A2(new_n286_), .A3(new_n613_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1331gat));
  NOR2_X1   g571(.A1(new_n452_), .A2(new_n471_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n699_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT110), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G57gat), .B1(new_n776_), .B2(new_n425_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n688_), .A2(new_n690_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n254_), .A3(new_n773_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n778_), .A2(KEYINPUT111), .A3(new_n254_), .A4(new_n773_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n425_), .A2(G57gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n777_), .B1(new_n783_), .B2(new_n784_), .ZN(G1332gat));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n700_), .A3(new_n782_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G64gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G64gat), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n581_), .A2(G64gat), .ZN(new_n790_));
  OAI22_X1  g589(.A1(new_n788_), .A2(new_n789_), .B1(new_n775_), .B2(new_n790_), .ZN(G1333gat));
  NAND3_X1  g590(.A1(new_n776_), .A2(new_n625_), .A3(new_n651_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n651_), .A3(new_n782_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(G71gat), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(G71gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(G1334gat));
  NAND3_X1  g596(.A1(new_n781_), .A2(new_n613_), .A3(new_n782_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G78gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G78gat), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n647_), .A2(G78gat), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n800_), .A2(new_n801_), .B1(new_n775_), .B2(new_n802_), .ZN(G1335gat));
  NAND2_X1  g602(.A1(new_n773_), .A2(new_n255_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n746_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(G85gat), .B1(new_n805_), .B2(new_n425_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT43), .B1(new_n686_), .B2(new_n736_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n678_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n424_), .A2(new_n315_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n806_), .B1(new_n809_), .B2(new_n810_), .ZN(G1336gat));
  AOI21_X1  g610(.A(G92gat), .B1(new_n805_), .B2(new_n700_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n581_), .A2(new_n316_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n809_), .B2(new_n813_), .ZN(G1337gat));
  OAI211_X1 g613(.A(new_n255_), .B(new_n773_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G99gat), .B1(new_n815_), .B2(new_n642_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n805_), .A2(new_n312_), .A3(new_n651_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n299_), .B1(new_n809_), .B2(new_n651_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n818_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT113), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n822_), .A3(KEYINPUT51), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n820_), .A2(new_n821_), .A3(KEYINPUT51), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n823_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n827_), .B2(new_n824_), .ZN(G1338gat));
  NAND3_X1  g627(.A1(new_n805_), .A2(new_n298_), .A3(new_n613_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n298_), .B1(new_n809_), .B2(new_n613_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n831_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1339gat));
  NAND2_X1  g635(.A1(new_n427_), .A2(new_n433_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n435_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT55), .A3(new_n434_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n434_), .A2(KEYINPUT55), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n443_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT56), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n837_), .B2(new_n435_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n445_), .B1(new_n844_), .B2(new_n434_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n840_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n842_), .A2(new_n847_), .A3(new_n471_), .A4(new_n446_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n235_), .A2(new_n297_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n297_), .B1(new_n220_), .B2(new_n229_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n457_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n235_), .A2(KEYINPUT79), .A3(new_n297_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n467_), .B1(new_n853_), .B2(new_n462_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n454_), .B(new_n462_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n461_), .A2(new_n455_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(KEYINPUT116), .A3(new_n467_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(new_n857_), .A3(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n860_), .A2(KEYINPUT117), .A3(new_n470_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT117), .B1(new_n860_), .B2(new_n470_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n447_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n848_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT57), .B1(new_n864_), .B2(new_n689_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866_));
  AOI211_X1 g665(.A(new_n866_), .B(new_n687_), .C1(new_n848_), .C2(new_n863_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  AND4_X1   g667(.A1(new_n846_), .A2(new_n839_), .A3(new_n840_), .A4(new_n443_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n846_), .B1(new_n845_), .B2(new_n840_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT116), .B1(new_n858_), .B2(new_n467_), .ZN(new_n873_));
  AOI211_X1 g672(.A(new_n855_), .B(new_n469_), .C1(new_n461_), .C2(new_n455_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n857_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n470_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n872_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n860_), .A2(KEYINPUT117), .A3(new_n470_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n871_), .A2(KEYINPUT58), .A3(new_n880_), .A4(new_n446_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884_));
  INV_X1    g683(.A(new_n880_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n842_), .A2(new_n446_), .A3(new_n847_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n886_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n888_), .A2(KEYINPUT118), .A3(KEYINPUT58), .A4(new_n880_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n883_), .A2(new_n737_), .A3(new_n887_), .A4(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n868_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n255_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n264_), .B1(new_n341_), .B2(new_n353_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n261_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n361_), .B1(new_n895_), .B2(new_n362_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n357_), .A2(new_n359_), .A3(KEYINPUT37), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n472_), .B(new_n254_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT54), .B1(new_n898_), .B2(new_n453_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n364_), .A2(new_n900_), .A3(new_n472_), .A4(new_n452_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n648_), .B1(new_n892_), .B2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n700_), .A2(new_n424_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G113gat), .B1(new_n906_), .B2(new_n471_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n905_), .A2(KEYINPUT119), .A3(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n905_), .B2(KEYINPUT119), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n472_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n907_), .B1(new_n911_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g711(.A(G120gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n452_), .B2(KEYINPUT60), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(KEYINPUT60), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(KEYINPUT120), .B2(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n906_), .B(new_n916_), .C1(KEYINPUT120), .C2(new_n914_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n452_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n913_), .ZN(G1341gat));
  AOI21_X1  g718(.A(G127gat), .B1(new_n906_), .B2(new_n254_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n255_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g721(.A(G134gat), .B1(new_n906_), .B2(new_n687_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n736_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g724(.A1(new_n892_), .A2(new_n902_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n651_), .A2(new_n647_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n926_), .A2(new_n904_), .A3(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n471_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g730(.A1(new_n928_), .A2(new_n452_), .ZN(new_n932_));
  XOR2_X1   g731(.A(KEYINPUT121), .B(G148gat), .Z(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1345gat));
  OR3_X1    g733(.A1(new_n928_), .A2(G155gat), .A3(new_n255_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n936_));
  OAI21_X1  g735(.A(G155gat), .B1(new_n928_), .B2(new_n255_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1346gat));
  INV_X1    g739(.A(G162gat), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n928_), .A2(new_n941_), .A3(new_n736_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n929_), .A2(new_n687_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n941_), .B2(new_n943_), .ZN(G1347gat));
  AOI21_X1  g743(.A(new_n254_), .B1(new_n868_), .B2(new_n890_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n899_), .A2(new_n901_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n647_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n581_), .A2(new_n425_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n651_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n472_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(KEYINPUT123), .ZN(new_n951_));
  OAI21_X1  g750(.A(G169gat), .B1(new_n947_), .B2(new_n951_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n952_), .A2(KEYINPUT62), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(KEYINPUT62), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n950_), .A2(new_n536_), .ZN(new_n955_));
  OAI22_X1  g754(.A1(new_n953_), .A2(new_n954_), .B1(new_n947_), .B2(new_n955_), .ZN(G1348gat));
  NAND2_X1  g755(.A1(new_n947_), .A2(KEYINPUT124), .ZN(new_n957_));
  INV_X1    g756(.A(new_n949_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n959_), .B(new_n647_), .C1(new_n945_), .C2(new_n946_), .ZN(new_n960_));
  AND2_X1   g759(.A1(new_n453_), .A2(G176gat), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n957_), .A2(new_n958_), .A3(new_n960_), .A4(new_n961_), .ZN(new_n962_));
  OAI211_X1 g761(.A(new_n643_), .B(new_n948_), .C1(new_n945_), .C2(new_n946_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n535_), .B1(new_n963_), .B2(new_n452_), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1349gat));
  NAND4_X1  g764(.A1(new_n957_), .A2(new_n254_), .A3(new_n958_), .A4(new_n960_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n966_), .A2(new_n517_), .ZN(new_n967_));
  INV_X1    g766(.A(new_n549_), .ZN(new_n968_));
  NAND4_X1  g767(.A1(new_n903_), .A2(new_n254_), .A3(new_n968_), .A4(new_n948_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n963_), .ZN(new_n972_));
  NAND4_X1  g771(.A1(new_n972_), .A2(KEYINPUT125), .A3(new_n254_), .A4(new_n968_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n971_), .A2(new_n973_), .ZN(new_n974_));
  OAI21_X1  g773(.A(KEYINPUT126), .B1(new_n967_), .B2(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n966_), .A2(new_n517_), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977_));
  NAND4_X1  g776(.A1(new_n976_), .A2(new_n977_), .A3(new_n971_), .A4(new_n973_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n975_), .A2(new_n978_), .ZN(G1350gat));
  OAI21_X1  g778(.A(G190gat), .B1(new_n963_), .B2(new_n736_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n687_), .A2(new_n550_), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n980_), .B1(new_n963_), .B2(new_n981_), .ZN(G1351gat));
  NAND3_X1  g781(.A1(new_n926_), .A2(new_n927_), .A3(new_n948_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n983_), .A2(new_n472_), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n984_), .B(new_n484_), .ZN(G1352gat));
  INV_X1    g784(.A(new_n983_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n986_), .A2(new_n453_), .A3(new_n482_), .ZN(new_n987_));
  OAI21_X1  g786(.A(G204gat), .B1(new_n983_), .B2(new_n452_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n987_), .A2(new_n988_), .ZN(new_n989_));
  MUX2_X1   g788(.A(new_n987_), .B(new_n989_), .S(KEYINPUT127), .Z(G1353gat));
  NOR2_X1   g789(.A1(new_n983_), .A2(new_n255_), .ZN(new_n991_));
  NOR2_X1   g790(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n992_));
  AND2_X1   g791(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n993_));
  OAI21_X1  g792(.A(new_n991_), .B1(new_n992_), .B2(new_n993_), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n994_), .B1(new_n991_), .B2(new_n992_), .ZN(G1354gat));
  INV_X1    g794(.A(G218gat), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n983_), .A2(new_n996_), .A3(new_n736_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n986_), .A2(new_n687_), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n997_), .B1(new_n996_), .B2(new_n998_), .ZN(G1355gat));
endmodule


