//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n584_, new_n585_, new_n586_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  AND3_X1   g003(.A1(new_n204_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n206_));
  INV_X1    g005(.A(new_n202_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT84), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n205_), .B1(new_n206_), .B2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n212_), .B(KEYINPUT80), .Z(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT22), .B(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(G176gat), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n211_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT82), .B1(new_n204_), .B2(KEYINPUT23), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n208_), .B2(new_n207_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n204_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT83), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n213_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  INV_X1    g028(.A(G190gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT26), .B1(new_n230_), .B2(KEYINPUT79), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(KEYINPUT26), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n229_), .B(new_n231_), .C1(new_n232_), .C2(KEYINPUT79), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n228_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n225_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n224_), .A2(KEYINPUT83), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n218_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G197gat), .B(G204gat), .Z(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(KEYINPUT21), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(KEYINPUT21), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G211gat), .B(G218gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n240_), .A2(new_n241_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n237_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G226gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT19), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n217_), .B1(new_n222_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT26), .B(G190gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n229_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n223_), .B1(new_n227_), .B2(new_n212_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n210_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT20), .B1(new_n255_), .B2(new_n244_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n245_), .A2(new_n248_), .A3(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT91), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n255_), .B2(new_n244_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n237_), .B2(new_n244_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n247_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(KEYINPUT91), .A3(new_n258_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT18), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  NOR2_X1   g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G1gat), .B(G29gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G57gat), .B(G85gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G155gat), .B(G162gat), .Z(new_n279_));
  NAND3_X1  g078(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT87), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT3), .ZN(new_n283_));
  INV_X1    g082(.A(G141gat), .ZN(new_n284_));
  INV_X1    g083(.A(G148gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n282_), .B(new_n286_), .C1(new_n287_), .C2(KEYINPUT2), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n279_), .B1(new_n281_), .B2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT88), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n279_), .A2(new_n291_), .ZN(new_n292_));
  AND3_X1   g091(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n287_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n289_), .A2(KEYINPUT88), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n290_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT92), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n290_), .A2(new_n296_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n297_), .A2(new_n298_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT86), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT92), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n301_), .B1(new_n309_), .B2(new_n300_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n278_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(KEYINPUT4), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT4), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n307_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n312_), .B1(new_n316_), .B2(new_n311_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n270_), .A2(new_n272_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n311_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT93), .ZN(new_n321_));
  INV_X1    g120(.A(new_n311_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(new_n310_), .B2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(KEYINPUT93), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n277_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT33), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n319_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n328_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n326_), .A2(KEYINPUT95), .A3(KEYINPUT33), .A4(new_n277_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n318_), .A2(new_n329_), .A3(new_n330_), .A4(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT96), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n324_), .A2(new_n278_), .A3(new_n325_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n324_), .A2(KEYINPUT96), .A3(new_n278_), .A4(new_n325_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n269_), .A2(KEYINPUT32), .ZN(new_n337_));
  INV_X1    g136(.A(new_n245_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n247_), .B1(new_n338_), .B2(new_n256_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n262_), .A2(new_n247_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n265_), .B2(new_n337_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n335_), .A2(new_n336_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n332_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT85), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT30), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n237_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n306_), .B(KEYINPUT31), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G15gat), .B(G43gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n350_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n302_), .A2(KEYINPUT29), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n360_), .B(KEYINPUT28), .Z(new_n361_));
  AOI22_X1  g160(.A1(new_n302_), .A2(KEYINPUT29), .B1(new_n242_), .B2(new_n243_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT90), .ZN(new_n365_));
  INV_X1    g164(.A(G228gat), .ZN(new_n366_));
  OR2_X1    g165(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n365_), .B(new_n369_), .Z(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n363_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n359_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n265_), .B(new_n269_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  INV_X1    g177(.A(new_n272_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n339_), .A2(new_n340_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n380_), .B2(new_n271_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n377_), .A2(new_n378_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n374_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n358_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n373_), .A3(new_n356_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n383_), .A2(new_n385_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n344_), .A2(new_n376_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G229gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT73), .B(G15gat), .ZN(new_n389_));
  INV_X1    g188(.A(G22gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(KEYINPUT74), .B(G1gat), .Z(new_n392_));
  INV_X1    g191(.A(G8gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT14), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G8gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G29gat), .B(G36gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G43gat), .B(G50gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(new_n399_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n388_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT15), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n403_), .B(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT77), .B1(new_n400_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n403_), .B(KEYINPUT15), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n399_), .A4(new_n398_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n388_), .B(KEYINPUT78), .Z(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n407_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G113gat), .B(G141gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G169gat), .B(G197gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  XOR2_X1   g220(.A(new_n418_), .B(new_n421_), .Z(new_n422_));
  NOR2_X1   g221(.A1(new_n387_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G231gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n400_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT11), .ZN(new_n427_));
  INV_X1    g226(.A(G57gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(G64gat), .ZN(new_n429_));
  INV_X1    g228(.A(G64gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(G57gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n427_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(G57gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(G64gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(KEYINPUT11), .ZN(new_n435_));
  XOR2_X1   g234(.A(G71gat), .B(G78gat), .Z(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G71gat), .B(G78gat), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n439_), .A2(KEYINPUT11), .A3(new_n433_), .A4(new_n434_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n437_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n438_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n426_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT76), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G127gat), .B(G155gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n446_), .B(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G183gat), .B(G211gat), .Z(new_n451_));
  AND2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n450_), .A2(new_n451_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n424_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n450_), .A2(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n451_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n445_), .A2(new_n424_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT7), .ZN(new_n460_));
  INV_X1    g259(.A(G99gat), .ZN(new_n461_));
  INV_X1    g260(.A(G106gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n468_), .A2(new_n470_), .A3(KEYINPUT64), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT64), .B1(new_n468_), .B2(new_n470_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n466_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G85gat), .B(G92gat), .Z(new_n474_));
  OR2_X1    g273(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n468_), .A2(new_n470_), .ZN(new_n479_));
  OAI211_X1 g278(.A(KEYINPUT66), .B(new_n474_), .C1(new_n479_), .C2(new_n465_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT8), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n468_), .A2(new_n470_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT66), .B1(new_n483_), .B2(new_n474_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n478_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n474_), .A2(KEYINPUT9), .ZN(new_n486_));
  INV_X1    g285(.A(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  OR3_X1    g287(.A1(new_n487_), .A2(new_n488_), .A3(KEYINPUT9), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT10), .B(G99gat), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n486_), .B(new_n489_), .C1(G106gat), .C2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n471_), .A2(new_n472_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n485_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n411_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT34), .ZN(new_n497_));
  OAI221_X1 g296(.A(new_n495_), .B1(KEYINPUT35), .B2(new_n497_), .C1(new_n405_), .C2(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(KEYINPUT35), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  XNOR2_X1  g299(.A(G190gat), .B(G218gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n500_), .A2(KEYINPUT36), .A3(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(KEYINPUT36), .Z(new_n505_));
  AND2_X1   g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT37), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n459_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT13), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n494_), .A2(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n443_), .A2(new_n485_), .A3(new_n493_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n437_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n442_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n485_), .A2(new_n493_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n516_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G230gat), .A2(G233gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT71), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT71), .ZN(new_n525_));
  INV_X1    g324(.A(new_n523_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n491_), .A2(new_n492_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n483_), .A2(new_n474_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(KEYINPUT8), .A3(new_n480_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n531_), .B2(new_n478_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n525_), .B(new_n526_), .C1(new_n532_), .C2(new_n443_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .A4(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n522_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT69), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT69), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n536_), .C1(new_n517_), .C2(new_n520_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G120gat), .B(G148gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT5), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G176gat), .B(G204gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(KEYINPUT72), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n542_), .A2(new_n549_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n514_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n552_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(KEYINPUT13), .A3(new_n550_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n513_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n423_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n335_), .A2(new_n336_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n559_), .A2(new_n561_), .A3(new_n392_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT97), .Z(new_n563_));
  INV_X1    g362(.A(KEYINPUT38), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n562_), .B(KEYINPUT97), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT38), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n344_), .A2(new_n376_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n386_), .A2(new_n382_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n507_), .B(KEYINPUT98), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n556_), .A2(new_n422_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n570_), .A2(new_n459_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(G1gat), .B1(new_n574_), .B2(new_n560_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n565_), .A2(new_n567_), .A3(new_n575_), .ZN(G1324gat));
  NOR3_X1   g375(.A1(new_n558_), .A2(G8gat), .A3(new_n382_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G8gat), .B1(new_n574_), .B2(new_n382_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(KEYINPUT39), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(KEYINPUT39), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n577_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(new_n582_), .Z(G1325gat));
  OAI21_X1  g382(.A(G15gat), .B1(new_n574_), .B2(new_n359_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT41), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n558_), .A2(G15gat), .A3(new_n359_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(G1326gat));
  OAI21_X1  g386(.A(G22gat), .B1(new_n574_), .B2(new_n374_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT42), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n559_), .A2(new_n390_), .A3(new_n373_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(G1327gat));
  INV_X1    g390(.A(new_n422_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n459_), .A2(new_n556_), .A3(new_n508_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n570_), .A2(KEYINPUT100), .A3(new_n592_), .A4(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n375_), .B1(new_n332_), .B2(new_n343_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n383_), .A2(new_n385_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n382_), .A2(new_n596_), .A3(new_n560_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n592_), .B(new_n593_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n594_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(G29gat), .B1(new_n601_), .B2(new_n561_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT43), .B1(new_n387_), .B2(new_n512_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT43), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n507_), .B(KEYINPUT37), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n604_), .B(new_n605_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n573_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n459_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT44), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611_));
  INV_X1    g410(.A(new_n609_), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n611_), .B(new_n612_), .C1(new_n603_), .C2(new_n606_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n561_), .A2(G29gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n602_), .B1(new_n614_), .B2(new_n615_), .ZN(G1328gat));
  NOR2_X1   g415(.A1(new_n382_), .A2(G36gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n594_), .A2(new_n600_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n594_), .A2(new_n600_), .A3(KEYINPUT102), .A4(new_n617_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n622_));
  AND3_X1   g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(G36gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n382_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n614_), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n625_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n620_), .A2(new_n621_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n622_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n610_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n613_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n627_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G36gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n629_), .B1(new_n636_), .B2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n631_), .A2(new_n641_), .ZN(G1329gat));
  INV_X1    g441(.A(new_n359_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G43gat), .B1(new_n601_), .B2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n643_), .A2(G43gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n614_), .B2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g446(.A(G50gat), .B1(new_n601_), .B2(new_n373_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n373_), .A2(G50gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n614_), .B2(new_n649_), .ZN(G1331gat));
  INV_X1    g449(.A(new_n556_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n592_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n570_), .A2(new_n459_), .A3(new_n572_), .A4(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G57gat), .B1(new_n653_), .B2(new_n560_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n387_), .A2(new_n592_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n458_), .A2(new_n454_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n556_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n561_), .A2(new_n428_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(G1332gat));
  OAI21_X1  g458(.A(G64gat), .B1(new_n653_), .B2(new_n382_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT48), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n627_), .A2(new_n430_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n661_), .B1(new_n657_), .B2(new_n662_), .ZN(G1333gat));
  OR3_X1    g462(.A1(new_n657_), .A2(G71gat), .A3(new_n359_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G71gat), .B1(new_n653_), .B2(new_n359_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT105), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n666_), .A2(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n664_), .B1(new_n669_), .B2(new_n670_), .ZN(G1334gat));
  OR3_X1    g470(.A1(new_n657_), .A2(G78gat), .A3(new_n374_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G78gat), .B1(new_n653_), .B2(new_n374_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT50), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n673_), .A2(KEYINPUT50), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT106), .ZN(G1335gat));
  INV_X1    g477(.A(new_n459_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n652_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT107), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n607_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G85gat), .B1(new_n682_), .B2(new_n560_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n459_), .A2(new_n651_), .A3(new_n508_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n655_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n487_), .A3(new_n561_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n687_), .ZN(G1336gat));
  OAI21_X1  g487(.A(G92gat), .B1(new_n682_), .B2(new_n382_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n686_), .A2(new_n488_), .A3(new_n627_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1337gat));
  OAI21_X1  g490(.A(G99gat), .B1(new_n682_), .B2(new_n359_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n359_), .A2(new_n490_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n685_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n462_), .A3(new_n373_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n607_), .A2(new_n681_), .A3(new_n373_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT52), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(G106gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n697_), .B2(G106gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g501(.A1(new_n627_), .A2(new_n560_), .A3(new_n383_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT114), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT55), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n534_), .B2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n521_), .A2(new_n533_), .A3(new_n524_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n709_), .B2(new_n536_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n710_), .B2(new_n535_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n521_), .A2(new_n533_), .A3(new_n524_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n712_), .A2(KEYINPUT109), .A3(KEYINPUT55), .A4(new_n522_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n546_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT56), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n713_), .B(new_n708_), .C1(new_n535_), .C2(new_n710_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(KEYINPUT56), .A3(new_n546_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n534_), .A2(new_n547_), .A3(new_n540_), .A4(new_n538_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n414_), .A2(new_n404_), .A3(new_n416_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n404_), .A2(new_n406_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n421_), .B1(new_n723_), .B2(new_n415_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n418_), .A2(new_n421_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n721_), .A2(new_n725_), .A3(KEYINPUT111), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT111), .B1(new_n721_), .B2(new_n725_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT58), .ZN(new_n731_));
  AOI22_X1  g530(.A1(new_n720_), .A2(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n731_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n733_), .B(new_n728_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n605_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT113), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n605_), .B(new_n737_), .C1(new_n732_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n592_), .A2(new_n721_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n718_), .A2(KEYINPUT56), .A3(new_n546_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT56), .B1(new_n718_), .B2(new_n546_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n725_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n507_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT57), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n740_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n745_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n508_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT57), .B1(new_n752_), .B2(KEYINPUT110), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n749_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n705_), .B1(new_n739_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n748_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(KEYINPUT110), .A3(KEYINPUT57), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n758_), .A2(KEYINPUT114), .A3(new_n736_), .A4(new_n738_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n679_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT54), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n557_), .A2(new_n422_), .A3(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n656_), .A2(new_n422_), .A3(new_n651_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n761_), .A2(KEYINPUT54), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n761_), .A2(KEYINPUT54), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n704_), .B1(new_n760_), .B2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G113gat), .B1(new_n769_), .B2(new_n592_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n760_), .A2(new_n768_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n703_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT59), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT59), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n763_), .A2(new_n767_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n459_), .B1(new_n758_), .B2(new_n735_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n774_), .B(new_n703_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n773_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n592_), .A2(G113gat), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT115), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n770_), .B1(new_n778_), .B2(new_n780_), .ZN(G1340gat));
  INV_X1    g580(.A(G120gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n651_), .B2(KEYINPUT60), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n769_), .B(new_n783_), .C1(KEYINPUT60), .C2(new_n782_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n778_), .A2(new_n556_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n786_), .B2(new_n782_), .ZN(G1341gat));
  OAI211_X1 g586(.A(new_n459_), .B(new_n777_), .C1(new_n769_), .C2(new_n774_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G127gat), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n772_), .A2(G127gat), .A3(new_n679_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n790_), .A3(KEYINPUT116), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1342gat));
  NAND2_X1  g594(.A1(new_n778_), .A2(new_n605_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(G134gat), .ZN(new_n797_));
  OR3_X1    g596(.A1(new_n772_), .A2(G134gat), .A3(new_n572_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1343gat));
  NAND3_X1  g598(.A1(new_n758_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n459_), .B1(new_n800_), .B2(new_n705_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n775_), .B1(new_n801_), .B2(new_n759_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n385_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n382_), .A3(new_n561_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n422_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(new_n284_), .ZN(G1344gat));
  NOR2_X1   g605(.A1(new_n804_), .A2(new_n651_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(new_n285_), .ZN(G1345gat));
  NOR2_X1   g607(.A1(new_n804_), .A2(new_n679_), .ZN(new_n809_));
  XOR2_X1   g608(.A(KEYINPUT61), .B(G155gat), .Z(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(G1346gat));
  INV_X1    g610(.A(G162gat), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n804_), .A2(new_n812_), .A3(new_n512_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n804_), .B2(new_n572_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT117), .B(new_n812_), .C1(new_n804_), .C2(new_n572_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(G1347gat));
  OR2_X1    g617(.A1(new_n775_), .A2(new_n776_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n561_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n592_), .A3(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n215_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(G169gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(KEYINPUT62), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(KEYINPUT62), .B2(new_n823_), .ZN(G1348gat));
  NOR2_X1   g624(.A1(new_n561_), .A2(new_n382_), .ZN(new_n826_));
  AND4_X1   g625(.A1(G176gat), .A2(new_n826_), .A3(new_n643_), .A4(new_n556_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n771_), .B2(new_n374_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT119), .B(new_n373_), .C1(new_n760_), .C2(new_n768_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT120), .B(new_n827_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n556_), .B(new_n820_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n832_));
  INV_X1    g631(.A(G176gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT118), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n836_), .A3(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT119), .B1(new_n802_), .B2(new_n373_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n771_), .A2(new_n828_), .A3(new_n374_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT120), .B1(new_n842_), .B2(new_n827_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT121), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n827_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n831_), .A4(new_n838_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n844_), .A2(new_n849_), .ZN(G1349gat));
  NAND2_X1  g649(.A1(new_n819_), .A2(new_n820_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n851_), .A2(new_n229_), .A3(new_n679_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n842_), .A2(new_n643_), .A3(new_n459_), .A4(new_n826_), .ZN(new_n853_));
  INV_X1    g652(.A(G183gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n851_), .B2(new_n512_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n571_), .A2(new_n251_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT122), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n851_), .B2(new_n858_), .ZN(G1351gat));
  AND2_X1   g658(.A1(new_n803_), .A2(new_n826_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n592_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n556_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT123), .B(G204gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1353gat));
  NOR2_X1   g664(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT124), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(KEYINPUT125), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n860_), .A2(new_n459_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(KEYINPUT125), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT126), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n870_), .B(new_n872_), .ZN(G1354gat));
  AOI21_X1  g672(.A(G218gat), .B1(new_n860_), .B2(new_n571_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n605_), .A2(G218gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT127), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n860_), .B2(new_n876_), .ZN(G1355gat));
endmodule


