//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT9), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT10), .ZN(new_n214_));
  INV_X1    g013(.A(G99gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n220_), .A3(new_n217_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT64), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n213_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT66), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT66), .B1(new_n203_), .B2(new_n205_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n215_), .A3(new_n220_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n225_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT65), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n209_), .A2(new_n235_), .A3(new_n210_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT8), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n237_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n230_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n206_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT8), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n239_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n224_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT11), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT67), .B(G71gat), .ZN(new_n247_));
  INV_X1    g046(.A(G78gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(G78gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n244_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G230gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT68), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n244_), .B2(new_n255_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n244_), .A2(new_n255_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n222_), .B(new_n219_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT69), .B1(new_n265_), .B2(new_n213_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n221_), .A2(new_n223_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n268_));
  INV_X1    g067(.A(new_n213_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n234_), .A2(new_n236_), .A3(new_n242_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n206_), .B2(new_n240_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n206_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT66), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n240_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n239_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n273_), .B1(new_n278_), .B2(KEYINPUT8), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n264_), .B1(new_n271_), .B2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n262_), .A2(new_n257_), .A3(new_n263_), .A4(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n282_));
  INV_X1    g081(.A(new_n263_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n244_), .A2(new_n255_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n282_), .B(new_n258_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G120gat), .B(G148gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT5), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G176gat), .B(G204gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n260_), .A2(new_n281_), .A3(new_n285_), .A4(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n281_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n282_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n289_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT13), .B1(new_n291_), .B2(new_n294_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT37), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G232gat), .A2(G233gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT34), .Z(new_n304_));
  XOR2_X1   g103(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G29gat), .B(G36gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G43gat), .B(G50gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT15), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n307_), .B(new_n308_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT15), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n266_), .A2(new_n270_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n238_), .A2(new_n243_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n224_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n242_), .B1(new_n277_), .B2(new_n239_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n318_), .B(new_n311_), .C1(new_n319_), .C2(new_n273_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n304_), .A2(new_n305_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n306_), .B1(new_n317_), .B2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n266_), .B(new_n270_), .C1(new_n319_), .C2(new_n273_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n306_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n321_), .A4(new_n320_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n302_), .B1(new_n323_), .B2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G190gat), .B(G218gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(G134gat), .B(G162gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT36), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n323_), .B2(new_n327_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(KEYINPUT36), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n328_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n335_), .ZN(new_n337_));
  AOI221_X4 g136(.A(new_n302_), .B1(new_n337_), .B2(new_n333_), .C1(new_n323_), .C2(new_n327_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n301_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n328_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n323_), .A2(new_n327_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n333_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n343_), .A3(new_n337_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n328_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(KEYINPUT37), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G127gat), .B(G155gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT16), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G183gat), .B(G211gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT72), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G15gat), .B(G22gat), .ZN(new_n354_));
  INV_X1    g153(.A(G1gat), .ZN(new_n355_));
  INV_X1    g154(.A(G8gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT14), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G1gat), .B(G8gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n353_), .B(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(G231gat), .A2(G233gat), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n254_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n255_), .A3(new_n364_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n351_), .A2(new_n352_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n347_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n300_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT73), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G183gat), .ZN(new_n376_));
  INV_X1    g175(.A(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n375_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G169gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(KEYINPUT81), .ZN(new_n383_));
  INV_X1    g182(.A(G169gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT81), .B1(new_n384_), .B2(KEYINPUT22), .ZN(new_n385_));
  INV_X1    g184(.A(G176gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n380_), .B(new_n381_), .C1(new_n383_), .C2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(KEYINPUT24), .A3(new_n381_), .A4(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n376_), .A2(KEYINPUT25), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G183gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n377_), .A2(KEYINPUT26), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT26), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G190gat), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n393_), .A2(new_n395_), .A3(new_n396_), .A4(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(new_n399_), .A3(KEYINPUT80), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n375_), .A2(new_n379_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n390_), .A2(new_n391_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT24), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT80), .B1(new_n392_), .B2(new_n399_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n388_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT84), .B(G197gat), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(G204gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G211gat), .B(G218gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT21), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n415_), .A2(new_n416_), .A3(G204gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n412_), .B1(G197gat), .B2(G204gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n411_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(G204gat), .B1(new_n415_), .B2(new_n416_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n408_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT21), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n414_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n414_), .B(KEYINPUT85), .C1(new_n420_), .C2(new_n423_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n407_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n380_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n375_), .A2(new_n378_), .A3(KEYINPUT88), .A4(new_n379_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n382_), .A2(new_n386_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n430_), .A2(new_n381_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n401_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n403_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n434_), .A2(new_n392_), .A3(new_n399_), .A4(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n424_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT20), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n428_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n424_), .B1(new_n437_), .B2(KEYINPUT95), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(KEYINPUT95), .B2(new_n437_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n426_), .A2(new_n407_), .A3(new_n427_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(KEYINPUT20), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n444_), .B2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G8gat), .B(G36gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G64gat), .B(G92gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n443_), .A2(KEYINPUT20), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n448_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n444_), .B1(new_n428_), .B2(new_n440_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n448_), .A3(KEYINPUT89), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n455_), .A4(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(KEYINPUT27), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n455_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT91), .A3(new_n464_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT27), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n462_), .A2(new_n463_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n455_), .A4(new_n461_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT96), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT96), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n470_), .A2(new_n477_), .A3(new_n471_), .A4(new_n474_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n466_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G127gat), .B(G134gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G113gat), .B(G120gat), .Z(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G113gat), .B(G120gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT82), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT2), .ZN(new_n487_));
  INV_X1    g286(.A(G141gat), .ZN(new_n488_));
  INV_X1    g287(.A(G148gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT3), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .A4(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G155gat), .A2(G162gat), .ZN(new_n496_));
  OR2_X1    g295(.A1(G155gat), .A2(G162gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G141gat), .B(G148gat), .Z(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(KEYINPUT1), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n497_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n496_), .A2(KEYINPUT1), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT82), .B1(new_n481_), .B2(new_n482_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n486_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n480_), .B(new_n484_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n503_), .A3(new_n498_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(KEYINPUT92), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n505_), .B1(new_n508_), .B2(KEYINPUT82), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n504_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G225gat), .A2(G233gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n507_), .A2(KEYINPUT4), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n522_), .B2(new_n515_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G29gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G85gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT0), .B(G57gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n523_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G227gat), .A2(G233gat), .ZN(new_n529_));
  INV_X1    g328(.A(G15gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT30), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G71gat), .B(G99gat), .ZN(new_n533_));
  INV_X1    g332(.A(G43gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n532_), .A2(new_n535_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(new_n407_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n511_), .B(KEYINPUT31), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT83), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n541_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n539_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n538_), .A2(new_n407_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n538_), .A2(new_n407_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G22gat), .B(G50gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n504_), .A2(KEYINPUT29), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n424_), .ZN(new_n553_));
  INV_X1    g352(.A(G228gat), .ZN(new_n554_));
  INV_X1    g353(.A(G233gat), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n426_), .A2(new_n427_), .A3(new_n552_), .A4(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT86), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n551_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n559_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT86), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n551_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n504_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT28), .B1(new_n504_), .B2(KEYINPUT29), .ZN(new_n570_));
  XOR2_X1   g369(.A(G78gat), .B(G106gat), .Z(new_n571_));
  AND3_X1   g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n571_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n563_), .A2(new_n568_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n563_), .B2(new_n568_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n550_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n563_), .A2(new_n568_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n574_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n575_), .A3(new_n549_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n528_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n470_), .A2(new_n474_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(KEYINPUT33), .ZN(new_n586_));
  INV_X1    g385(.A(new_n521_), .ZN(new_n587_));
  AND4_X1   g386(.A1(new_n512_), .A2(new_n486_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n512_), .B1(new_n511_), .B2(new_n504_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n509_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n587_), .B1(new_n590_), .B2(new_n519_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n517_), .B1(new_n591_), .B2(new_n516_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n527_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n586_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n527_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n522_), .B2(new_n515_), .ZN(new_n597_));
  NOR4_X1   g396(.A1(new_n520_), .A2(KEYINPUT94), .A3(new_n516_), .A4(new_n521_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n595_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n586_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n523_), .A2(new_n527_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n523_), .B(new_n593_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n455_), .A2(KEYINPUT32), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n472_), .A2(new_n461_), .A3(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n450_), .B2(new_n604_), .ZN(new_n606_));
  OAI22_X1  g405(.A1(new_n584_), .A2(new_n602_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n581_), .A2(new_n575_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n550_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n479_), .A2(new_n583_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n310_), .A2(new_n360_), .A3(new_n313_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n358_), .A2(new_n359_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n358_), .A2(new_n359_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n311_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n612_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n360_), .A2(new_n309_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n616_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT74), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(KEYINPUT74), .A3(new_n616_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n613_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n617_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(G113gat), .B(G141gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(G169gat), .B(G197gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT77), .B1(new_n625_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n622_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT74), .B1(new_n618_), .B2(new_n616_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n624_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n612_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT77), .ZN(new_n637_));
  INV_X1    g436(.A(new_n630_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(new_n635_), .A3(new_n630_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT78), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT78), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n634_), .A2(new_n642_), .A3(new_n635_), .A4(new_n630_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n631_), .A2(new_n639_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n611_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n372_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n355_), .A3(new_n528_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n631_), .A2(new_n639_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n641_), .A2(new_n643_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n299_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT97), .ZN(new_n654_));
  INV_X1    g453(.A(new_n369_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n336_), .A2(new_n657_), .A3(new_n338_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT98), .B1(new_n344_), .B2(new_n345_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n611_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n656_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n603_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n647_), .A2(new_n648_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n649_), .A2(new_n665_), .A3(new_n666_), .ZN(G1324gat));
  INV_X1    g466(.A(new_n479_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n646_), .A2(new_n356_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n670_));
  OAI21_X1  g469(.A(G8gat), .B1(new_n670_), .B2(KEYINPUT99), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n663_), .B2(new_n668_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n672_), .A2(KEYINPUT99), .A3(new_n670_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(KEYINPUT99), .B2(new_n670_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n669_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(KEYINPUT40), .B(new_n669_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n664_), .B2(new_n549_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n646_), .A2(new_n530_), .A3(new_n550_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(G22gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n646_), .A2(new_n686_), .A3(new_n609_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n663_), .A2(new_n609_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(G22gat), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G22gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1327gat));
  NOR2_X1   g493(.A1(new_n654_), .A2(new_n369_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n611_), .B2(new_n347_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n476_), .A2(new_n478_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n465_), .A3(new_n583_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n607_), .A2(new_n610_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  INV_X1    g500(.A(new_n347_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n696_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n695_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707_), .B2(new_n603_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n300_), .A2(new_n660_), .A3(new_n369_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n645_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n603_), .A2(G29gat), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT103), .Z(new_n713_));
  OAI21_X1  g512(.A(new_n708_), .B1(new_n711_), .B2(new_n713_), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n711_), .A2(G36gat), .A3(new_n479_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT45), .Z(new_n716_));
  OAI21_X1  g515(.A(G36gat), .B1(new_n707_), .B2(new_n479_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(KEYINPUT46), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  OAI21_X1  g521(.A(new_n534_), .B1(new_n711_), .B2(new_n549_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n550_), .A2(G43gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n707_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g525(.A1(new_n711_), .A2(G50gat), .A3(new_n608_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n707_), .A2(new_n608_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G50gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n728_), .A2(new_n729_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(G1331gat));
  NAND4_X1  g532(.A1(new_n662_), .A2(new_n644_), .A3(new_n300_), .A4(new_n369_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT106), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(G57gat), .A3(new_n528_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n737_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n370_), .A2(new_n299_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n741_), .A2(KEYINPUT105), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n611_), .A2(new_n652_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(KEYINPUT105), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G57gat), .B1(new_n746_), .B2(new_n528_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n738_), .A2(new_n739_), .A3(new_n747_), .ZN(G1332gat));
  NAND2_X1  g547(.A1(new_n735_), .A2(new_n668_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G64gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  OR3_X1    g551(.A1(new_n745_), .A2(G64gat), .A3(new_n479_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1333gat));
  INV_X1    g553(.A(G71gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n735_), .B2(new_n550_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n550_), .A2(new_n755_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT110), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n745_), .B2(new_n760_), .ZN(G1334gat));
  AOI21_X1  g560(.A(new_n248_), .B1(new_n735_), .B2(new_n609_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n746_), .A2(new_n248_), .A3(new_n609_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1335gat));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n300_), .A2(new_n644_), .A3(new_n655_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n704_), .B2(new_n769_), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT112), .B(new_n768_), .C1(new_n696_), .C2(new_n703_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n603_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n299_), .A2(new_n660_), .A3(new_n369_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n743_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n207_), .A3(new_n528_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1336gat));
  OAI21_X1  g576(.A(G92gat), .B1(new_n772_), .B2(new_n479_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n208_), .A3(new_n668_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1337gat));
  NAND3_X1  g579(.A1(new_n775_), .A2(new_n550_), .A3(new_n218_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n550_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G99gat), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT51), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT113), .B(new_n782_), .C1(new_n783_), .C2(G99gat), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n701_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT43), .B(new_n347_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n769_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT112), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n704_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n549_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n790_), .B(new_n781_), .C1(new_n796_), .C2(new_n215_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n787_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n781_), .B1(new_n796_), .B2(new_n215_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n790_), .B1(new_n799_), .B2(KEYINPUT113), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n784_), .A2(new_n785_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n798_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n789_), .A2(new_n802_), .ZN(G1338gat));
  NAND3_X1  g602(.A1(new_n775_), .A2(new_n220_), .A3(new_n609_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G106gat), .B1(new_n793_), .B2(new_n608_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(KEYINPUT52), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(KEYINPUT52), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n804_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n652_), .A2(new_n291_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n281_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n281_), .B2(new_n812_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n324_), .A2(new_n264_), .B1(new_n244_), .B2(new_n255_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n257_), .B1(new_n816_), .B2(new_n262_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n814_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n811_), .B1(new_n818_), .B2(new_n290_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n281_), .A2(new_n812_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT55), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n281_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n817_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n289_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n810_), .B1(new_n819_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n612_), .A2(new_n616_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n613_), .B1(new_n827_), .B2(KEYINPUT116), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(KEYINPUT116), .B2(new_n827_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n630_), .B1(new_n623_), .B2(new_n613_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n641_), .A2(new_n643_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n295_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT57), .B(new_n660_), .C1(new_n826_), .C2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n660_), .B1(new_n826_), .B2(new_n833_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n292_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n644_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n817_), .B1(new_n820_), .B2(KEYINPUT55), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n811_), .B(new_n290_), .C1(new_n842_), .C2(new_n822_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT56), .B1(new_n824_), .B2(new_n289_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n832_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n660_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n831_), .A2(new_n291_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT58), .B(new_n848_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n702_), .A3(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n836_), .A2(new_n839_), .A3(new_n847_), .A4(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n655_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n299_), .A2(new_n347_), .A3(new_n644_), .A4(new_n369_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n578_), .A2(new_n603_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n860_), .A2(new_n479_), .A3(new_n861_), .A4(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n858_), .B1(new_n854_), .B2(new_n655_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n861_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n864_), .A2(new_n668_), .A3(new_n865_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n867_));
  OAI21_X1  g666(.A(new_n863_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n644_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n866_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n860_), .A2(new_n479_), .A3(new_n861_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT118), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n644_), .A2(G113gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n869_), .B1(new_n874_), .B2(new_n875_), .ZN(G1340gat));
  OAI211_X1 g675(.A(new_n863_), .B(new_n300_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G120gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n299_), .A2(KEYINPUT60), .ZN(new_n879_));
  INV_X1    g678(.A(G120gat), .ZN(new_n880_));
  MUX2_X1   g679(.A(KEYINPUT60), .B(new_n879_), .S(new_n880_), .Z(new_n881_));
  NAND3_X1  g680(.A1(new_n871_), .A2(new_n873_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT120), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n878_), .A2(new_n885_), .A3(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1341gat));
  OAI21_X1  g686(.A(G127gat), .B1(new_n868_), .B2(new_n655_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n655_), .A2(G127gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n874_), .B2(new_n889_), .ZN(G1342gat));
  OAI21_X1  g689(.A(G134gat), .B1(new_n868_), .B2(new_n347_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n660_), .A2(G134gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n874_), .B2(new_n892_), .ZN(G1343gat));
  NOR4_X1   g692(.A1(new_n864_), .A2(new_n668_), .A3(new_n603_), .A4(new_n582_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n652_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT121), .B(G141gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n300_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g698(.A1(new_n894_), .A2(new_n369_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n894_), .A2(new_n903_), .A3(new_n661_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n894_), .A2(new_n702_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1347gat));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n479_), .A2(new_n528_), .A3(new_n578_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n860_), .A2(new_n652_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n860_), .A2(KEYINPUT122), .A3(new_n652_), .A4(new_n908_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n911_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n908_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n864_), .A2(new_n644_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n382_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n384_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n918_));
  AOI21_X1  g717(.A(KEYINPUT62), .B1(new_n918_), .B2(new_n912_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n907_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n921_));
  OAI21_X1  g720(.A(G169gat), .B1(new_n915_), .B2(KEYINPUT122), .ZN(new_n922_));
  INV_X1    g721(.A(new_n912_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n924_), .A2(KEYINPUT123), .A3(new_n916_), .A4(new_n913_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n920_), .A2(new_n925_), .ZN(G1348gat));
  NOR2_X1   g725(.A1(new_n864_), .A2(new_n914_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n300_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G176gat), .ZN(G1349gat));
  NOR3_X1   g728(.A1(new_n864_), .A2(new_n655_), .A3(new_n914_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(G183gat), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n393_), .A2(new_n395_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n930_), .ZN(G1350gat));
  AOI21_X1  g732(.A(new_n377_), .B1(new_n927_), .B2(new_n702_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT124), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n927_), .A2(new_n396_), .A3(new_n398_), .A4(new_n661_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n582_), .A2(new_n528_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT125), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n864_), .A2(new_n479_), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n652_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n300_), .ZN(new_n943_));
  XOR2_X1   g742(.A(KEYINPUT126), .B(G204gat), .Z(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1353gat));
  AND2_X1   g744(.A1(new_n940_), .A2(new_n369_), .ZN(new_n946_));
  XOR2_X1   g745(.A(KEYINPUT63), .B(G211gat), .Z(new_n947_));
  AOI21_X1  g746(.A(KEYINPUT127), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n947_), .ZN(new_n949_));
  OR2_X1    g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n946_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n948_), .B1(new_n951_), .B2(KEYINPUT127), .ZN(G1354gat));
  INV_X1    g751(.A(G218gat), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n940_), .A2(new_n953_), .A3(new_n661_), .ZN(new_n954_));
  AND2_X1   g753(.A1(new_n940_), .A2(new_n702_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n955_), .B2(new_n953_), .ZN(G1355gat));
endmodule


