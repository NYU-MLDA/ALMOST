//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT18), .B(G64gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT20), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT96), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n218_), .A2(new_n219_), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT24), .B1(new_n214_), .B2(new_n215_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT96), .B1(new_n227_), .B2(new_n224_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n216_), .A2(new_n217_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n230_), .A2(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n231_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT97), .ZN(new_n241_));
  NAND2_X1  g040(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT97), .B1(new_n244_), .B2(new_n239_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n238_), .B1(new_n246_), .B2(new_n213_), .ZN(new_n247_));
  INV_X1    g046(.A(G183gat), .ZN(new_n248_));
  INV_X1    g047(.A(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n222_), .A2(new_n223_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT98), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n235_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  INV_X1    g055(.A(G204gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G197gat), .ZN(new_n258_));
  INV_X1    g057(.A(G197gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G204gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n258_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n259_), .A2(G204gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n263_), .B2(KEYINPUT90), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT90), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n260_), .A3(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n256_), .B(new_n262_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n256_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT21), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n210_), .B1(new_n255_), .B2(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n270_), .A2(new_n272_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n218_), .A2(KEYINPUT81), .A3(new_n225_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n227_), .B2(new_n224_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n237_), .A2(KEYINPUT24), .A3(new_n214_), .A4(new_n215_), .ZN(new_n279_));
  OR3_X1    g078(.A1(new_n249_), .A2(KEYINPUT78), .A3(KEYINPUT26), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT26), .B1(new_n249_), .B2(KEYINPUT78), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n232_), .A3(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n276_), .A2(new_n278_), .A3(new_n279_), .A4(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n213_), .B1(new_n244_), .B2(new_n239_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(new_n237_), .A3(new_n251_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n275_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n209_), .B1(new_n274_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n285_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n273_), .A2(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n235_), .A2(new_n254_), .A3(new_n270_), .A4(new_n272_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT20), .A4(new_n209_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n206_), .B1(new_n287_), .B2(new_n292_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n229_), .A2(new_n234_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT20), .B1(new_n275_), .B2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n273_), .A2(new_n288_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n208_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n206_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(new_n291_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT27), .B1(new_n293_), .B2(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n287_), .A2(new_n292_), .A3(new_n206_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT20), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n208_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT102), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n274_), .A2(new_n286_), .A3(new_n209_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT102), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n306_), .A3(new_n208_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n301_), .B1(new_n308_), .B2(new_n206_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n300_), .B1(new_n309_), .B2(KEYINPUT27), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT93), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G228gat), .A2(G233gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(KEYINPUT92), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(KEYINPUT86), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  AND4_X1   g123(.A1(new_n319_), .A2(new_n320_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n326_), .A2(KEYINPUT85), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT85), .B1(new_n326_), .B2(new_n327_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n316_), .B1(new_n325_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n332_));
  INV_X1    g131(.A(G155gat), .ZN(new_n333_));
  INV_X1    g132(.A(G162gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n338_), .A3(new_n336_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT84), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT84), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n335_), .A2(new_n338_), .A3(new_n342_), .A4(new_n336_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n326_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n346_), .A2(new_n347_), .B1(G141gat), .B2(G148gat), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n331_), .A2(new_n337_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n273_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n313_), .A2(KEYINPUT92), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n314_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n314_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n344_), .A2(new_n348_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT85), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n319_), .A2(new_n320_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n315_), .B(new_n337_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n354_), .B1(new_n361_), .B2(new_n273_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n312_), .B1(new_n353_), .B2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G78gat), .B(G106gat), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n351_), .A2(new_n314_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n361_), .A2(new_n273_), .B1(KEYINPUT92), .B2(new_n313_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT93), .B(new_n366_), .C1(new_n367_), .C2(new_n314_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT94), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n371_));
  XOR2_X1   g170(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G22gat), .B(G50gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n349_), .A2(new_n350_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n355_), .A2(new_n350_), .A3(new_n359_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n374_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n373_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n378_), .A3(new_n373_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n371_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n371_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n383_), .A2(new_n379_), .A3(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT94), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n363_), .A2(new_n368_), .A3(new_n387_), .A4(new_n365_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n364_), .B(new_n366_), .C1(new_n367_), .C2(new_n314_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT95), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n353_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n392_), .A2(KEYINPUT95), .A3(new_n364_), .A4(new_n366_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n370_), .A2(new_n386_), .A3(new_n388_), .A4(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n365_), .B1(new_n353_), .B2(new_n362_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n389_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n385_), .B2(new_n382_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n311_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G127gat), .B(G134gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n360_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n355_), .A2(new_n359_), .A3(new_n403_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(KEYINPUT4), .A3(new_n406_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n408_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n360_), .A2(new_n412_), .A3(new_n404_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G1gat), .B(G29gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT100), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n415_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n409_), .A2(new_n414_), .A3(new_n421_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT103), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT103), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n409_), .A2(new_n414_), .A3(new_n426_), .A4(new_n421_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n425_), .A2(KEYINPUT104), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT104), .B1(new_n425_), .B2(new_n427_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G71gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n403_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT30), .B(G99gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G15gat), .B(G43gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT31), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n288_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n436_), .B(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n400_), .A2(new_n430_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n425_), .A2(KEYINPUT104), .A3(new_n427_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n425_), .A2(new_n427_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT104), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n399_), .A2(new_n442_), .A3(new_n445_), .A4(new_n310_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT105), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n424_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT101), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(KEYINPUT33), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n293_), .A2(new_n299_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n424_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n410_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n407_), .A2(new_n411_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n422_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n451_), .A2(new_n452_), .A3(new_n454_), .A4(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n450_), .B1(new_n449_), .B2(KEYINPUT33), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n298_), .A2(KEYINPUT32), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n308_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n425_), .A2(new_n461_), .A3(new_n427_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n287_), .A2(new_n292_), .A3(new_n460_), .ZN(new_n463_));
  OAI22_X1  g262(.A1(new_n458_), .A2(new_n459_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n399_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n430_), .A2(KEYINPUT105), .A3(new_n399_), .A4(new_n310_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n448_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n440_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n441_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G57gat), .B(G64gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT11), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G71gat), .B(G78gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT11), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n471_), .B(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n476_), .B2(new_n473_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G85gat), .B(G92gat), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT9), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT6), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT10), .B(G99gat), .Z(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT9), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(G85gat), .A3(G92gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n482_), .A2(KEYINPUT64), .A3(new_n485_), .A4(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT64), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n479_), .A2(new_n487_), .A3(new_n481_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n485_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  OR3_X1    g293(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n481_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n478_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n496_), .B2(new_n478_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n477_), .B1(new_n493_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G230gat), .A2(G233gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(new_n478_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT8), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n496_), .A2(new_n497_), .A3(new_n478_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n477_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n488_), .A4(new_n492_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n488_), .A3(new_n492_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT12), .A3(new_n477_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n503_), .A2(new_n504_), .A3(new_n510_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT65), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n510_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n501_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n513_), .B1(new_n517_), .B2(new_n504_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G120gat), .B(G148gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT67), .ZN(new_n520_));
  XOR2_X1   g319(.A(G176gat), .B(G204gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n518_), .A2(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n513_), .B(new_n524_), .C1(new_n517_), .C2(new_n504_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT13), .Z(new_n529_));
  XNOR2_X1  g328(.A(G190gat), .B(G218gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G43gat), .B(G50gat), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(G36gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537_));
  INV_X1    g336(.A(G36gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT69), .B(G29gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n536_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n541_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n545_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n511_), .A2(new_n547_), .A3(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n548_), .A2(new_n549_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n508_), .A2(new_n559_), .A3(new_n488_), .A4(new_n492_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n551_), .A2(KEYINPUT71), .A3(new_n558_), .A4(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n493_), .A2(new_n500_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n550_), .A2(new_n547_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n560_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(new_n565_), .B2(new_n556_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n551_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n534_), .B(new_n561_), .C1(new_n566_), .C2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT72), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n555_), .B1(new_n551_), .B2(new_n560_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n567_), .B1(new_n571_), .B2(new_n562_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n534_), .A4(new_n561_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n534_), .B1(new_n572_), .B2(new_n561_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n533_), .B2(new_n532_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(new_n577_), .A3(KEYINPUT37), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G15gat), .B(G22gat), .ZN(new_n583_));
  INV_X1    g382(.A(G1gat), .ZN(new_n584_));
  INV_X1    g383(.A(G8gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT14), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G1gat), .B(G8gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n477_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(G211gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(KEYINPUT16), .B(G183gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT73), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n596_), .A2(new_n597_), .ZN(new_n602_));
  OR3_X1    g401(.A1(new_n592_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT74), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n582_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G169gat), .B(G197gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT77), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n589_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n589_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT75), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n550_), .A2(new_n547_), .A3(new_n589_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT76), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n550_), .A2(new_n547_), .A3(KEYINPUT76), .A4(new_n589_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n625_), .A2(new_n618_), .A3(new_n615_), .A4(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(new_n620_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n613_), .B(new_n622_), .C1(new_n628_), .C2(new_n621_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n621_), .B1(new_n627_), .B2(new_n620_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n622_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n612_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR4_X1   g433(.A1(new_n470_), .A2(new_n529_), .A3(new_n608_), .A4(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n430_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n584_), .A3(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT38), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n529_), .A2(new_n634_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n604_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n468_), .A2(new_n469_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n441_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n642_), .B1(new_n645_), .B2(new_n578_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n578_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n470_), .A2(KEYINPUT106), .A3(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n641_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT107), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n642_), .A3(new_n578_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT106), .B1(new_n470_), .B2(new_n647_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(KEYINPUT107), .A3(new_n641_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n430_), .B1(new_n651_), .B2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n638_), .B1(new_n656_), .B2(new_n584_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT108), .Z(G1324gat));
  OAI21_X1  g457(.A(G8gat), .B1(new_n649_), .B2(new_n310_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT39), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n635_), .A2(new_n585_), .A3(new_n311_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1325gat));
  AOI21_X1  g463(.A(KEYINPUT107), .B1(new_n654_), .B2(new_n641_), .ZN(new_n665_));
  AOI211_X1 g464(.A(new_n650_), .B(new_n640_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n440_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G15gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G15gat), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G15gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n635_), .A2(new_n673_), .A3(new_n440_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n674_), .A3(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n635_), .A2(new_n677_), .A3(new_n399_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n465_), .B1(new_n651_), .B2(new_n655_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n679_), .A2(KEYINPUT42), .A3(new_n677_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n399_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(G22gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n680_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT111), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n686_), .B(new_n678_), .C1(new_n680_), .C2(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n645_), .A2(new_n582_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(KEYINPUT43), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(KEYINPUT43), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n639_), .B(new_n606_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n689_), .B(KEYINPUT43), .ZN(new_n696_));
  INV_X1    g495(.A(new_n694_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n696_), .A2(new_n639_), .A3(new_n606_), .A4(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n636_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT113), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT113), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n695_), .A2(new_n698_), .A3(new_n701_), .A4(new_n636_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(G29gat), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n606_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n470_), .A2(new_n578_), .A3(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n639_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n430_), .A2(G29gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n703_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NAND3_X1  g508(.A1(new_n695_), .A2(new_n311_), .A3(new_n698_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n310_), .B(KEYINPUT114), .Z(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n538_), .A3(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT45), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n711_), .A2(KEYINPUT46), .A3(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  NAND4_X1  g518(.A1(new_n695_), .A2(new_n698_), .A3(G43gat), .A4(new_n440_), .ZN(new_n720_));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n707_), .B2(new_n469_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1330gat));
  NAND3_X1  g524(.A1(new_n695_), .A2(new_n399_), .A3(new_n698_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G50gat), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n707_), .A2(G50gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n465_), .B2(new_n728_), .ZN(G1331gat));
  INV_X1    g528(.A(new_n529_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n608_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT116), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n634_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n470_), .B(new_n733_), .C1(new_n732_), .C2(new_n731_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n636_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n730_), .A2(new_n633_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n654_), .A2(new_n704_), .A3(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n636_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n735_), .B1(G57gat), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n740_), .A3(new_n712_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n712_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G64gat), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT48), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT48), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1333gat));
  NAND3_X1  g545(.A1(new_n734_), .A2(new_n431_), .A3(new_n440_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n737_), .A2(new_n440_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(G71gat), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT49), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT49), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n734_), .A2(new_n753_), .A3(new_n399_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n737_), .A2(new_n399_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(G78gat), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT50), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT50), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  AND2_X1   g558(.A1(new_n705_), .A2(new_n736_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n636_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n696_), .A2(new_n606_), .A3(new_n736_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n636_), .A2(G85gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n760_), .B2(new_n311_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n762_), .A2(new_n203_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(new_n712_), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n762_), .B2(new_n469_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(new_n440_), .A3(new_n483_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n760_), .A2(new_n484_), .A3(new_n399_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n696_), .A2(new_n399_), .A3(new_n606_), .A4(new_n736_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G106gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  NAND3_X1  g581(.A1(new_n607_), .A2(new_n730_), .A3(new_n634_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n625_), .A2(new_n615_), .A3(new_n626_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n619_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n615_), .A2(new_n618_), .A3(new_n616_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n611_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n630_), .A2(new_n631_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(new_n611_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n503_), .A2(new_n512_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT55), .A3(new_n504_), .A4(new_n510_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n504_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n503_), .A2(new_n512_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n515_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n513_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n525_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n525_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n527_), .B(new_n791_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n582_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n804_), .B2(new_n582_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n802_), .A2(new_n803_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n528_), .A2(new_n791_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n633_), .A2(KEYINPUT117), .A3(new_n527_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT117), .B1(new_n633_), .B2(new_n527_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n800_), .A2(new_n801_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n810_), .B1(new_n818_), .B2(new_n647_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n815_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n813_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n800_), .A2(new_n801_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n811_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n578_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n809_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n604_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n785_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n400_), .A2(new_n636_), .A3(new_n440_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830_), .B2(new_n633_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n606_), .B1(new_n809_), .B2(new_n825_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n785_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT119), .B(new_n606_), .C1(new_n809_), .C2(new_n825_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  INV_X1    g637(.A(new_n829_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT59), .B1(new_n828_), .B2(new_n829_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(new_n633_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n831_), .B1(new_n843_), .B2(G113gat), .ZN(G1340gat));
  NAND3_X1  g643(.A1(new_n840_), .A2(new_n529_), .A3(new_n841_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT120), .B(G120gat), .Z(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n846_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n730_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n830_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT121), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n847_), .A2(new_n853_), .A3(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n830_), .B2(new_n704_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n842_), .A2(G127gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n604_), .ZN(G1342gat));
  AOI21_X1  g657(.A(G134gat), .B1(new_n830_), .B2(new_n647_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n582_), .A2(G134gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT122), .Z(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n842_), .B2(new_n861_), .ZN(G1343gat));
  NOR3_X1   g661(.A1(new_n828_), .A2(new_n465_), .A3(new_n712_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n430_), .A2(new_n440_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n633_), .A3(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT123), .B(G141gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1344gat));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n529_), .A3(new_n864_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT124), .B(G148gat), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n868_), .B(new_n869_), .Z(G1345gat));
  NAND3_X1  g669(.A1(new_n863_), .A2(new_n704_), .A3(new_n864_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  AND4_X1   g672(.A1(G162gat), .A2(new_n863_), .A3(new_n582_), .A4(new_n864_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n863_), .A2(new_n647_), .A3(new_n864_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n334_), .B2(new_n875_), .ZN(G1347gat));
  INV_X1    g675(.A(new_n712_), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n877_), .A2(new_n636_), .A3(new_n399_), .A4(new_n469_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n837_), .A2(new_n633_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G169gat), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n880_), .A2(KEYINPUT62), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(KEYINPUT62), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n837_), .A2(KEYINPUT125), .A3(new_n878_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT125), .B1(new_n837_), .B2(new_n878_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n633_), .A2(new_n246_), .ZN(new_n886_));
  OAI22_X1  g685(.A1(new_n881_), .A2(new_n882_), .B1(new_n885_), .B2(new_n886_), .ZN(G1348gat));
  INV_X1    g686(.A(new_n828_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n878_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n889_), .A2(new_n213_), .A3(new_n730_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n529_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n213_), .ZN(G1349gat));
  NOR2_X1   g691(.A1(new_n827_), .A2(new_n232_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n248_), .B1(new_n889_), .B2(new_n606_), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT126), .B(new_n893_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(G1350gat));
  INV_X1    g698(.A(new_n582_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G190gat), .B1(new_n885_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n647_), .A2(new_n233_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n885_), .B2(new_n902_), .ZN(G1351gat));
  NOR3_X1   g702(.A1(new_n828_), .A2(new_n440_), .A3(new_n877_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n636_), .A2(new_n465_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n634_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n259_), .ZN(G1352gat));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n730_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n257_), .ZN(G1353gat));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n906_), .A2(new_n827_), .A3(new_n911_), .A4(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n906_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n604_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n915_), .B2(new_n911_), .ZN(G1354gat));
  OAI21_X1  g715(.A(KEYINPUT127), .B1(new_n906_), .B2(new_n578_), .ZN(new_n917_));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n904_), .A2(new_n919_), .A3(new_n905_), .A4(new_n647_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n918_), .A3(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n914_), .A2(G218gat), .A3(new_n582_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1355gat));
endmodule


