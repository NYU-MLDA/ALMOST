//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  INV_X1    g002(.A(G50gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT69), .B(G43gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT15), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT10), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT10), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G99gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(G106gat), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT9), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  INV_X1    g023(.A(G92gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(KEYINPUT64), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n228_), .A3(KEYINPUT9), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n219_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n209_), .A3(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n233_), .A2(new_n216_), .A3(new_n217_), .A4(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n220_), .A2(new_n221_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT8), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n235_), .B(new_n236_), .C1(new_n238_), .C2(KEYINPUT8), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n230_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n208_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G232gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT34), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT35), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n230_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n207_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n246_), .A2(new_n247_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n251_), .B(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G190gat), .B(G218gat), .Z(new_n255_));
  XNOR2_X1  g054(.A(G134gat), .B(G162gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT71), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n254_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n257_), .B(KEYINPUT36), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n254_), .A2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n202_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n261_), .B(KEYINPUT37), .C1(new_n254_), .C2(new_n264_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G127gat), .B(G155gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(G211gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT16), .B(G183gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n273_));
  INV_X1    g072(.A(G57gat), .ZN(new_n274_));
  INV_X1    g073(.A(G64gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G57gat), .A2(G64gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281_));
  INV_X1    g080(.A(G78gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G71gat), .ZN(new_n283_));
  INV_X1    g082(.A(G71gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G78gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n280_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(new_n280_), .B2(new_n286_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n279_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n280_), .A2(new_n286_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT66), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n280_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n278_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G15gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G22gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT73), .B(G1gat), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G8gat), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n298_), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT74), .B1(new_n298_), .B2(KEYINPUT14), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n296_), .B(new_n302_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n305_));
  INV_X1    g104(.A(G231gat), .ZN(new_n306_));
  INV_X1    g105(.A(G233gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n309_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n294_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n294_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n310_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n272_), .B1(new_n317_), .B2(KEYINPUT17), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n272_), .A2(KEYINPUT17), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT75), .B1(new_n313_), .B2(new_n316_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI211_X1 g121(.A(KEYINPUT75), .B(KEYINPUT76), .C1(new_n313_), .C2(new_n316_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n318_), .B(new_n319_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n320_), .A2(new_n321_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n323_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT17), .B1(new_n313_), .B2(new_n316_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n272_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n319_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n326_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n268_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT77), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT23), .ZN(new_n335_));
  INV_X1    g134(.A(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT24), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(KEYINPUT24), .A3(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n335_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(KEYINPUT78), .B(G190gat), .Z(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(new_n344_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n342_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n335_), .B1(G183gat), .B2(new_n347_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351_));
  OR3_X1    g150(.A1(new_n351_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT80), .B(G176gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(G169gat), .B1(new_n351_), .B2(KEYINPUT79), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n340_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n349_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT30), .Z(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G15gat), .B(G43gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n359_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n358_), .B(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(new_n363_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT82), .B1(new_n365_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n363_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n360_), .A2(new_n364_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G134gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT81), .B(G127gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  INV_X1    g177(.A(G134gat), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n374_), .A2(new_n379_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n378_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT31), .Z(new_n384_));
  NAND3_X1  g183(.A1(new_n369_), .A2(new_n373_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  OAI211_X1 g185(.A(KEYINPUT82), .B(new_n386_), .C1(new_n365_), .C2(new_n368_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT86), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT21), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G197gat), .B(G204gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n390_), .A2(new_n394_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n396_), .B(new_n398_), .C1(KEYINPUT21), .C2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(KEYINPUT21), .A3(new_n397_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n405_));
  NAND3_X1  g204(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT1), .B1(new_n408_), .B2(new_n403_), .ZN(new_n409_));
  OR2_X1    g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n413_), .B(KEYINPUT3), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n412_), .B(KEYINPUT2), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n404_), .A2(new_n406_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n410_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT29), .ZN(new_n422_));
  NOR2_X1   g221(.A1(KEYINPUT85), .A2(G228gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(KEYINPUT85), .A2(G228gat), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n307_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n402_), .A2(new_n422_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n427_), .B1(new_n402_), .B2(new_n422_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G78gat), .B(G106gat), .Z(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G22gat), .B(G50gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n421_), .B2(KEYINPUT29), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n421_), .A2(KEYINPUT29), .A3(new_n436_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n435_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n439_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n431_), .B(new_n432_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n402_), .A2(new_n422_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n426_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n428_), .A3(new_n432_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n448_), .A2(KEYINPUT88), .A3(new_n442_), .A4(new_n440_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n433_), .B1(new_n445_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT89), .B1(new_n431_), .B2(new_n432_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n452_));
  INV_X1    g251(.A(new_n432_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n452_), .B(new_n453_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n450_), .B1(new_n443_), .B2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n415_), .A2(new_n377_), .A3(new_n420_), .A4(new_n382_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n415_), .A2(new_n420_), .B1(new_n377_), .B2(new_n382_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n421_), .A2(new_n383_), .A3(KEYINPUT91), .ZN(new_n462_));
  OAI211_X1 g261(.A(KEYINPUT92), .B(KEYINPUT4), .C1(new_n461_), .C2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466_));
  INV_X1    g265(.A(new_n462_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n421_), .A2(new_n383_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n458_), .A3(new_n457_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(new_n468_), .B2(KEYINPUT4), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n463_), .B(new_n465_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G57gat), .B(G85gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(G1gat), .B(G29gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n467_), .A2(new_n469_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n464_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT95), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n479_), .B1(new_n473_), .B2(new_n482_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n473_), .A2(new_n482_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(KEYINPUT95), .A3(new_n478_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n456_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G8gat), .B(G36gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(new_n225_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT18), .B(G64gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  NOR2_X1   g294(.A1(new_n402_), .A2(new_n357_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n344_), .A2(G190gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n343_), .A2(new_n345_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n342_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n335_), .B1(G183gat), .B2(G190gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT22), .B(G169gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n353_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n340_), .A3(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n496_), .A2(new_n497_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G226gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT19), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT90), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n402_), .A2(new_n357_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n400_), .A2(new_n505_), .A3(new_n401_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT20), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n514_), .A2(new_n516_), .A3(new_n509_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n495_), .B1(new_n512_), .B2(new_n517_), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n514_), .A2(new_n516_), .A3(new_n509_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n495_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n519_), .B(new_n520_), .C1(new_n511_), .C2(new_n507_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT27), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n518_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT94), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n516_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n515_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n513_), .A3(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n528_), .A2(new_n509_), .B1(new_n511_), .B2(new_n507_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n524_), .B1(new_n529_), .B2(new_n520_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n513_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT94), .B1(new_n515_), .B2(KEYINPUT20), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n509_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n507_), .A2(new_n511_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(KEYINPUT96), .A3(new_n495_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n521_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n523_), .B1(new_n537_), .B2(KEYINPUT27), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n491_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n488_), .A2(new_n478_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n484_), .A3(new_n483_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n520_), .A2(KEYINPUT32), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  OR3_X1    g342(.A1(new_n512_), .A2(new_n542_), .A3(new_n517_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n541_), .A2(new_n489_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n518_), .A2(new_n521_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n463_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n464_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n548_), .B(new_n479_), .C1(new_n464_), .C2(new_n481_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT33), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n486_), .A2(new_n550_), .ZN(new_n551_));
  AOI211_X1 g350(.A(KEYINPUT33), .B(new_n479_), .C1(new_n473_), .C2(new_n482_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n546_), .B(new_n549_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n456_), .B1(new_n545_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n388_), .B1(new_n539_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n487_), .A2(new_n490_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n388_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n456_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n537_), .A2(KEYINPUT27), .ZN(new_n559_));
  INV_X1    g358(.A(new_n523_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n555_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n333_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n249_), .A2(new_n294_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n242_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(KEYINPUT12), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n315_), .A2(new_n568_), .A3(new_n242_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n565_), .A2(new_n566_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n571_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT68), .ZN(new_n578_));
  XOR2_X1   g377(.A(G176gat), .B(G204gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n572_), .A2(new_n575_), .A3(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n304_), .A2(new_n305_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(new_n207_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(G229gat), .A3(G233gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n208_), .A2(new_n305_), .A3(new_n304_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n207_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G169gat), .B(G197gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n598_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n587_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n564_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n556_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n297_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n262_), .A2(new_n265_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT97), .B1(new_n563_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n331_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n563_), .A2(KEYINPUT97), .A3(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n602_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n556_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(G1gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n606_), .A2(new_n607_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n608_), .A2(new_n618_), .A3(new_n619_), .ZN(G1324gat));
  INV_X1    g419(.A(new_n602_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n613_), .A2(new_n621_), .A3(new_n538_), .A4(new_n614_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(new_n623_), .A3(G8gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n622_), .B2(G8gat), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n561_), .A2(G8gat), .ZN(new_n626_));
  OAI22_X1  g425(.A1(new_n624_), .A2(new_n625_), .B1(new_n604_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI221_X1 g428(.A(KEYINPUT40), .B1(new_n604_), .B2(new_n626_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1325gat));
  INV_X1    g430(.A(G15gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n388_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n603_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n616_), .B2(new_n633_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n636_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(G1326gat));
  INV_X1    g438(.A(G22gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n603_), .A2(new_n640_), .A3(new_n456_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n616_), .A2(new_n456_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(G22gat), .ZN(new_n644_));
  AOI211_X1 g443(.A(KEYINPUT42), .B(new_n640_), .C1(new_n616_), .C2(new_n456_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n644_), .B2(new_n645_), .ZN(G1327gat));
  AOI21_X1  g445(.A(new_n610_), .B1(new_n555_), .B2(new_n562_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n602_), .A2(new_n331_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n556_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n266_), .A2(new_n267_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n555_), .B2(new_n562_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n268_), .A2(KEYINPUT99), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n652_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n563_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n655_), .B1(new_n660_), .B2(KEYINPUT43), .ZN(new_n661_));
  INV_X1    g460(.A(new_n648_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n651_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n654_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n561_), .A2(new_n605_), .A3(new_n456_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n545_), .A2(new_n553_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n558_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n633_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n561_), .A2(new_n558_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(new_n556_), .A3(new_n388_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n664_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n555_), .A2(new_n562_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n653_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(KEYINPUT44), .A3(new_n648_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n663_), .A2(G29gat), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n650_), .B1(new_n675_), .B2(new_n556_), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n663_), .A2(new_n538_), .A3(new_n674_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n647_), .A2(new_n679_), .A3(new_n648_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n680_), .A2(KEYINPUT100), .A3(new_n561_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT100), .B1(new_n680_), .B2(new_n561_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(KEYINPUT45), .A3(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n682_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n678_), .A2(new_n683_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n678_), .A2(KEYINPUT46), .A3(new_n686_), .A4(new_n683_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1329gat));
  XOR2_X1   g490(.A(KEYINPUT101), .B(G43gat), .Z(new_n692_));
  INV_X1    g491(.A(new_n649_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n388_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n663_), .A2(new_n674_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n633_), .A2(G43gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g497(.A1(new_n649_), .A2(new_n204_), .A3(new_n456_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n663_), .A2(new_n456_), .A3(new_n674_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(G50gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n700_), .B2(G50gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1331gat));
  NOR2_X1   g503(.A1(new_n587_), .A2(new_n601_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n564_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n274_), .B1(new_n708_), .B2(new_n605_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  NOR4_X1   g511(.A1(new_n615_), .A2(new_n274_), .A3(new_n605_), .A4(new_n706_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(G1332gat));
  NAND3_X1  g513(.A1(new_n707_), .A2(new_n275_), .A3(new_n538_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n615_), .A2(new_n706_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n538_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(G64gat), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT48), .B(new_n275_), .C1(new_n717_), .C2(new_n538_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n715_), .B1(new_n719_), .B2(new_n720_), .ZN(G1333gat));
  NAND4_X1  g520(.A1(new_n613_), .A2(new_n633_), .A3(new_n614_), .A4(new_n705_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n722_), .A2(new_n723_), .A3(G71gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n722_), .B2(G71gat), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n707_), .A2(new_n284_), .A3(new_n633_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n726_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(G1334gat));
  NAND3_X1  g529(.A1(new_n707_), .A2(new_n282_), .A3(new_n456_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT50), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n717_), .A2(new_n456_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G78gat), .ZN(new_n734_));
  AOI211_X1 g533(.A(KEYINPUT50), .B(new_n282_), .C1(new_n717_), .C2(new_n456_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1335gat));
  NOR2_X1   g535(.A1(new_n706_), .A2(new_n331_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n647_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n556_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n661_), .A2(KEYINPUT106), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n661_), .A2(KEYINPUT106), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n737_), .A3(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(new_n224_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n741_), .B1(new_n745_), .B2(new_n556_), .ZN(G1336gat));
  AOI21_X1  g545(.A(G92gat), .B1(new_n740_), .B2(new_n538_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n744_), .A2(new_n225_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n538_), .ZN(G1337gat));
  NAND4_X1  g548(.A1(new_n742_), .A2(new_n633_), .A3(new_n737_), .A4(new_n743_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G99gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n210_), .A2(new_n212_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n740_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n633_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT108), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n751_), .A2(new_n754_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(KEYINPUT107), .A2(KEYINPUT51), .ZN(new_n758_));
  AOI22_X1  g557(.A1(G99gat), .A2(new_n750_), .B1(new_n753_), .B2(new_n633_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(KEYINPUT108), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n757_), .A2(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(G1338gat));
  NOR3_X1   g560(.A1(new_n706_), .A2(new_n558_), .A3(new_n331_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n653_), .B1(new_n563_), .B2(new_n659_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT109), .B(new_n762_), .C1(new_n763_), .C2(new_n655_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT109), .B1(new_n673_), .B2(new_n762_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n767_), .A2(G106gat), .A3(new_n770_), .A4(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n740_), .A2(new_n232_), .A3(new_n456_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774_));
  INV_X1    g573(.A(new_n762_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n661_), .B2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(G106gat), .A3(new_n771_), .A4(new_n764_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n769_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n772_), .A2(new_n773_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n772_), .A2(new_n778_), .A3(new_n773_), .A4(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  NOR3_X1   g582(.A1(new_n669_), .A2(new_n605_), .A3(new_n388_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n574_), .A2(KEYINPUT113), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n570_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n567_), .A2(new_n569_), .A3(new_n786_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n571_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n572_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n574_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT112), .B1(new_n795_), .B2(KEYINPUT55), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n792_), .A2(new_n794_), .A3(KEYINPUT114), .A4(new_n796_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n583_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT56), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n799_), .A2(new_n803_), .A3(new_n583_), .A4(new_n800_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n802_), .A2(new_n601_), .A3(new_n585_), .A4(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n589_), .A2(new_n592_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n591_), .A2(new_n593_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n806_), .B(new_n598_), .C1(new_n592_), .C2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n599_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n586_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n805_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n610_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n610_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n609_), .B1(new_n805_), .B2(new_n810_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n819_), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n585_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n801_), .B2(KEYINPUT56), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n809_), .A3(new_n804_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n823_), .A2(KEYINPUT58), .A3(new_n809_), .A4(new_n804_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n652_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT116), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n826_), .A2(new_n830_), .A3(new_n652_), .A4(new_n827_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n818_), .A2(new_n821_), .A3(new_n829_), .A4(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n612_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n599_), .A2(new_n600_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n331_), .A2(new_n834_), .A3(new_n587_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT111), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n331_), .A2(new_n834_), .A3(new_n837_), .A4(new_n587_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n268_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n785_), .B1(new_n833_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n601_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n832_), .B2(new_n612_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT59), .B1(new_n845_), .B2(new_n785_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n817_), .A2(new_n812_), .A3(new_n828_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n848_), .A2(new_n612_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n847_), .B(new_n784_), .C1(new_n849_), .C2(new_n841_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n846_), .A2(new_n601_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n844_), .B1(new_n851_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g651(.A(new_n587_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n853_), .B(new_n850_), .C1(new_n843_), .C2(new_n847_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n846_), .A2(KEYINPUT117), .A3(new_n853_), .A4(new_n850_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(G120gat), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n843_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(G1341gat));
  NOR3_X1   g661(.A1(new_n845_), .A2(new_n612_), .A3(new_n785_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864_));
  OR3_X1    g663(.A1(new_n863_), .A2(new_n864_), .A3(G127gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n863_), .B2(G127gat), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n846_), .A2(G127gat), .A3(new_n331_), .A4(new_n850_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(G1342gat));
  NOR3_X1   g667(.A1(new_n845_), .A2(new_n610_), .A3(new_n785_), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n869_), .A2(KEYINPUT119), .A3(G134gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT119), .B1(new_n869_), .B2(G134gat), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n846_), .A2(G134gat), .A3(new_n652_), .A4(new_n850_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(G1343gat));
  NOR3_X1   g672(.A1(new_n633_), .A2(new_n605_), .A3(new_n558_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT115), .B1(new_n819_), .B2(KEYINPUT57), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n820_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n829_), .A2(new_n831_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n331_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n561_), .B(new_n874_), .C1(new_n880_), .C2(new_n841_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n834_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT120), .B(G141gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n881_), .A2(new_n587_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT121), .B(G148gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1345gat));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n881_), .B2(new_n612_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n845_), .A2(new_n538_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n889_), .A2(new_n890_), .A3(new_n331_), .A4(new_n874_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n888_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1346gat));
  INV_X1    g694(.A(new_n881_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G162gat), .B1(new_n896_), .B2(new_n609_), .ZN(new_n897_));
  INV_X1    g696(.A(G162gat), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n896_), .B2(new_n899_), .ZN(G1347gat));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n841_), .B1(new_n612_), .B2(new_n848_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n557_), .A2(new_n538_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n456_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n903_), .A2(new_n834_), .A3(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n901_), .B(new_n902_), .C1(new_n907_), .C2(new_n336_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n502_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n601_), .B(new_n905_), .C1(new_n849_), .C2(new_n841_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n901_), .A2(new_n902_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n910_), .A2(G169gat), .A3(new_n911_), .A4(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n908_), .A2(new_n909_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT124), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n908_), .A2(new_n916_), .A3(new_n909_), .A4(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1348gat));
  OAI21_X1  g717(.A(new_n905_), .B1(new_n849_), .B2(new_n841_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n353_), .B1(new_n919_), .B2(new_n587_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n921_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n904_), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n845_), .A2(new_n337_), .A3(new_n587_), .A4(new_n456_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n922_), .A2(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(G1349gat));
  NOR3_X1   g725(.A1(new_n919_), .A2(new_n343_), .A3(new_n612_), .ZN(new_n927_));
  OR4_X1    g726(.A1(new_n456_), .A2(new_n845_), .A3(new_n612_), .A4(new_n904_), .ZN(new_n928_));
  INV_X1    g727(.A(G183gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n919_), .B2(new_n268_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n609_), .A2(new_n345_), .A3(new_n498_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n919_), .B2(new_n932_), .ZN(G1351gat));
  NOR2_X1   g732(.A1(new_n633_), .A2(new_n491_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n561_), .B1(new_n934_), .B2(KEYINPUT126), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n935_), .B(new_n937_), .C1(new_n880_), .C2(new_n841_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n834_), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n587_), .ZN(new_n941_));
  XOR2_X1   g740(.A(new_n941_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g741(.A1(new_n938_), .A2(new_n612_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(new_n943_), .B2(new_n944_), .ZN(G1354gat));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n948_), .B1(new_n938_), .B2(new_n610_), .ZN(new_n949_));
  INV_X1    g748(.A(G218gat), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n845_), .A2(new_n936_), .ZN(new_n951_));
  NAND4_X1  g750(.A1(new_n951_), .A2(KEYINPUT127), .A3(new_n609_), .A4(new_n935_), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n949_), .A2(new_n950_), .A3(new_n952_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n938_), .A2(new_n950_), .A3(new_n268_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1355gat));
endmodule


