//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT67), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n203_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n205_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n206_), .A2(new_n210_), .A3(KEYINPUT15), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(KEYINPUT9), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT6), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT6), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n221_), .A2(KEYINPUT9), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n219_), .A2(new_n222_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n220_), .A2(new_n221_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AOI211_X1 g033(.A(KEYINPUT8), .B(new_n230_), .C1(new_n234_), .C2(new_n227_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT7), .ZN(new_n237_));
  INV_X1    g036(.A(G99gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n217_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n225_), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n223_), .A2(KEYINPUT6), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n231_), .B(new_n239_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n230_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n236_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n229_), .B1(new_n235_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n215_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT34), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT35), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n229_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n224_), .A2(new_n226_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n239_), .A2(new_n231_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n243_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT8), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n242_), .A2(new_n236_), .A3(new_n243_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n206_), .A3(new_n210_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n246_), .A2(new_n251_), .A3(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n249_), .A2(new_n250_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n246_), .A2(new_n263_), .A3(new_n251_), .A4(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G190gat), .B(G218gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G134gat), .B(G162gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(KEYINPUT36), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n268_), .A2(KEYINPUT36), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n262_), .A2(new_n271_), .A3(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT27), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT76), .B(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT22), .B(G169gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G183gat), .ZN(new_n281_));
  INV_X1    g080(.A(G190gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT23), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(G183gat), .A3(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n282_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n280_), .A2(KEYINPUT89), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n276_), .A2(new_n277_), .B1(G169gat), .B2(G176gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT25), .B(G183gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G190gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G169gat), .ZN(new_n295_));
  INV_X1    g094(.A(G176gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n279_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n294_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  MUX2_X1   g099(.A(new_n286_), .B(new_n285_), .S(KEYINPUT78), .Z(new_n301_));
  AOI22_X1  g100(.A1(new_n288_), .A2(new_n291_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT21), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n304_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n308_), .A3(new_n306_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT90), .B1(new_n302_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n301_), .A2(new_n300_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n291_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n286_), .A2(new_n287_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n312_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT90), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n307_), .A2(new_n309_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n311_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n280_), .A2(KEYINPUT77), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n284_), .A2(KEYINPUT78), .A3(G183gat), .A4(G190gat), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(new_n287_), .C1(new_n286_), .C2(KEYINPUT78), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n289_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n300_), .A2(new_n286_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(KEYINPUT79), .A3(new_n327_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n310_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n320_), .A2(new_n332_), .A3(KEYINPUT20), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT18), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  NAND2_X1  g139(.A1(new_n330_), .A2(new_n331_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n318_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT91), .B1(new_n316_), .B2(new_n318_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT91), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n302_), .A2(new_n344_), .A3(new_n310_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n335_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n342_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n336_), .A2(new_n340_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n340_), .B1(new_n336_), .B2(new_n349_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n275_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G225gat), .A2(G233gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT3), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(G141gat), .B2(G148gat), .ZN(new_n360_));
  AND2_X1   g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n358_), .A2(new_n360_), .B1(KEYINPUT2), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT86), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT86), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G127gat), .B(G134gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT81), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n375_), .A2(new_n376_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n370_), .A2(KEYINPUT1), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n380_), .A2(KEYINPUT84), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(KEYINPUT84), .ZN(new_n382_));
  OAI221_X1 g181(.A(new_n369_), .B1(KEYINPUT1), .B2(new_n370_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n361_), .A2(new_n357_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n373_), .A2(new_n379_), .A3(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n375_), .B(new_n376_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n371_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n383_), .A2(new_n384_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n390_), .A3(KEYINPUT4), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n387_), .B(new_n392_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n353_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(G1gat), .B(G29gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT92), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n353_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n395_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n400_), .B1(new_n394_), .B2(new_n403_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n340_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n335_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n341_), .B2(new_n318_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n302_), .A2(KEYINPUT96), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n302_), .A2(KEYINPUT96), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n310_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  AND4_X1   g215(.A1(KEYINPUT20), .A2(new_n320_), .A3(new_n410_), .A4(new_n332_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n409_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n336_), .A2(new_n340_), .A3(new_n349_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT27), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n352_), .A2(new_n408_), .A3(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n388_), .A2(new_n389_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n318_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G228gat), .ZN(new_n425_));
  INV_X1    g224(.A(G233gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT87), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(KEYINPUT87), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n429_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n422_), .A2(new_n423_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT28), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n422_), .A2(new_n437_), .A3(new_n423_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n439_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n438_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n437_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n434_), .A2(KEYINPUT88), .A3(new_n440_), .A4(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n442_), .A2(new_n443_), .A3(new_n441_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n439_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n429_), .B(new_n432_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n444_), .A2(KEYINPUT88), .A3(new_n440_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n445_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n421_), .A2(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(KEYINPUT32), .B(new_n340_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n340_), .A2(KEYINPUT32), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n336_), .A2(new_n349_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n407_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT93), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n406_), .A2(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(KEYINPUT93), .B(new_n400_), .C1(new_n394_), .C2(new_n403_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n326_), .A2(KEYINPUT79), .A3(new_n327_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT79), .B1(new_n326_), .B2(new_n327_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n347_), .B1(new_n467_), .B2(new_n310_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n410_), .B1(new_n468_), .B2(new_n320_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n342_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n409_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT33), .B(new_n400_), .C1(new_n394_), .C2(new_n403_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n391_), .A2(new_n353_), .A3(new_n393_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n386_), .A2(new_n402_), .A3(new_n390_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n401_), .A3(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n471_), .A2(new_n472_), .A3(new_n419_), .A4(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n453_), .B(new_n459_), .C1(new_n464_), .C2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(G15gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n481_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n330_), .A2(new_n331_), .A3(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G71gat), .B(G99gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G43gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n482_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n478_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n482_), .A2(new_n484_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n488_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n482_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(KEYINPUT82), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n379_), .B(KEYINPUT31), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n491_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n478_), .B(new_n497_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n499_), .A2(KEYINPUT83), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT83), .B1(new_n499_), .B2(new_n500_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n455_), .A2(new_n477_), .A3(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n352_), .A2(new_n420_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n499_), .A2(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n505_), .A2(new_n408_), .A3(new_n453_), .A4(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n274_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G127gat), .B(G155gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT16), .ZN(new_n511_));
  XOR2_X1   g310(.A(G183gat), .B(G211gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G57gat), .B(G64gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT11), .ZN(new_n517_));
  XOR2_X1   g316(.A(G71gat), .B(G78gat), .Z(new_n518_));
  OR2_X1    g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n516_), .A2(KEYINPUT11), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n518_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G231gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528_));
  INV_X1    g327(.A(G8gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n527_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n524_), .B(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n533_), .A2(new_n514_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n515_), .B1(new_n534_), .B2(new_n513_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n535_), .B(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(new_n531_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n527_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n527_), .A2(new_n539_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n206_), .B(new_n210_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n215_), .B2(new_n532_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n532_), .A2(new_n211_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n542_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT72), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(KEYINPUT72), .A3(new_n548_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n545_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G113gat), .B(G141gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G169gat), .B(G197gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT65), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n521_), .A2(new_n520_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n517_), .A2(new_n518_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT66), .B1(new_n245_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT65), .B1(new_n245_), .B2(new_n565_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n562_), .A2(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT64), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n258_), .A2(new_n522_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT66), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n258_), .B2(new_n522_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(KEYINPUT65), .A3(KEYINPUT12), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n569_), .A2(new_n572_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n573_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n258_), .A2(new_n522_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n571_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G120gat), .B(G148gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT5), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n585_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND4_X1   g391(.A1(new_n509_), .A2(new_n538_), .A3(new_n561_), .A4(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n202_), .B1(new_n593_), .B2(new_n407_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT98), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n561_), .B(KEYINPUT75), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n535_), .B(new_n537_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n270_), .A2(new_n599_), .A3(new_n272_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT69), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n270_), .A2(new_n272_), .A3(new_n602_), .A4(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n269_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT68), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n272_), .B1(new_n606_), .B2(KEYINPUT68), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n598_), .B1(new_n604_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n597_), .A2(new_n592_), .A3(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT97), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n408_), .A2(G1gat), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n595_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT99), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n595_), .B(new_n620_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(G1324gat));
  XNOR2_X1  g421(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n623_));
  INV_X1    g422(.A(new_n505_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n593_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G8gat), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT39), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(KEYINPUT39), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n613_), .A2(new_n529_), .A3(new_n624_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n623_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n630_), .B(new_n623_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1325gat));
  INV_X1    g433(.A(new_n503_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n593_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G15gat), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n612_), .A2(G15gat), .A3(new_n503_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT101), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n453_), .B(KEYINPUT102), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n593_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n643_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n612_), .B2(new_n647_), .ZN(G1327gat));
  NAND2_X1  g447(.A1(new_n598_), .A2(new_n274_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT105), .Z(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(new_n592_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(new_n597_), .ZN(new_n652_));
  INV_X1    g451(.A(G29gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n407_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n604_), .A2(new_n610_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n592_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n561_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n659_), .A2(new_n538_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT44), .B1(new_n662_), .B2(KEYINPUT103), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n658_), .A2(new_n664_), .A3(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n658_), .A2(KEYINPUT44), .A3(new_n661_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n408_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n666_), .A2(new_n667_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G29gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n667_), .B1(new_n666_), .B2(new_n670_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n654_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n668_), .A2(new_n624_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n666_), .B2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n651_), .A2(new_n676_), .A3(new_n624_), .A4(new_n597_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n675_), .B1(new_n679_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n682_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n677_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n684_), .B(KEYINPUT46), .C1(new_n685_), .C2(new_n676_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1329gat));
  NAND2_X1  g486(.A1(new_n507_), .A2(G43gat), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n688_), .B(new_n669_), .C1(new_n663_), .C2(new_n665_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n652_), .A2(new_n635_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT107), .B(G43gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT47), .B1(new_n689_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n692_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n666_), .A2(new_n668_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n694_), .B(new_n695_), .C1(new_n696_), .C2(new_n688_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n693_), .A2(new_n697_), .ZN(G1330gat));
  AOI21_X1  g497(.A(G50gat), .B1(new_n652_), .B2(new_n644_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n696_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n454_), .A2(G50gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(G1331gat));
  INV_X1    g501(.A(new_n596_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n703_), .A2(new_n598_), .A3(new_n592_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n509_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n408_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n561_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n708_), .A2(new_n659_), .A3(new_n611_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n407_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n713_), .A3(new_n624_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G64gat), .B1(new_n706_), .B2(new_n505_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n716_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT109), .ZN(G1333gat));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n705_), .B2(new_n635_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT49), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n709_), .A2(new_n721_), .A3(new_n635_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1334gat));
  INV_X1    g524(.A(G78gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n705_), .B2(new_n644_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n709_), .A2(new_n726_), .A3(new_n644_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1335gat));
  AND2_X1   g529(.A1(new_n650_), .A2(new_n659_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(new_n708_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n407_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n733_), .A2(KEYINPUT110), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(KEYINPUT110), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n538_), .A2(new_n592_), .A3(new_n561_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n658_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT111), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n407_), .A2(G85gat), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT112), .Z(new_n740_));
  AOI22_X1  g539(.A1(new_n734_), .A2(new_n735_), .B1(new_n738_), .B2(new_n740_), .ZN(G1336gat));
  INV_X1    g540(.A(G92gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n732_), .A2(new_n742_), .A3(new_n624_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n738_), .A2(new_n624_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n742_), .ZN(G1337gat));
  AND3_X1   g544(.A1(new_n507_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n731_), .A2(new_n708_), .A3(new_n746_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT113), .Z(new_n748_));
  OAI21_X1  g547(.A(G99gat), .B1(new_n737_), .B2(new_n503_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT51), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n752_), .A3(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1338gat));
  NAND2_X1  g553(.A1(new_n504_), .A2(new_n508_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n606_), .A2(KEYINPUT68), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n607_), .A3(new_n272_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(KEYINPUT37), .A2(new_n757_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n657_), .B1(new_n755_), .B2(new_n758_), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT43), .B(new_n655_), .C1(new_n504_), .C2(new_n508_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n454_), .B(new_n736_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G106gat), .B1(new_n761_), .B2(new_n762_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n658_), .A2(KEYINPUT114), .A3(new_n454_), .A4(new_n736_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n762_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .A4(G106gat), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n732_), .A2(new_n217_), .A3(new_n454_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n774_), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  NAND3_X1  g575(.A1(new_n611_), .A2(new_n592_), .A3(new_n596_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n777_), .B(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n576_), .A2(new_n573_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n562_), .B1(new_n258_), .B2(new_n522_), .ZN(new_n782_));
  AOI22_X1  g581(.A1(KEYINPUT65), .A2(new_n575_), .B1(new_n782_), .B2(KEYINPUT12), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n571_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n569_), .A2(new_n573_), .A3(new_n576_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n571_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n577_), .A2(KEYINPUT55), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n566_), .A2(new_n562_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n578_), .B1(new_n790_), .B2(KEYINPUT12), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n572_), .A4(new_n569_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n785_), .A2(new_n788_), .B1(new_n789_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n780_), .B1(new_n794_), .B2(new_n585_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n585_), .A2(new_n780_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT116), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n786_), .A2(new_n787_), .A3(new_n571_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n787_), .B1(new_n786_), .B2(new_n571_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n789_), .A2(new_n793_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n799_), .B(new_n796_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n795_), .A2(new_n798_), .A3(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n660_), .A2(new_n587_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n215_), .A2(new_n532_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n542_), .A2(new_n548_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n558_), .B1(new_n547_), .B2(new_n543_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT117), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n813_), .B(new_n816_), .C1(new_n587_), .C2(new_n589_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n807_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n273_), .A2(KEYINPUT57), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n818_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n274_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n796_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n795_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n813_), .A2(new_n586_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n828_), .A2(KEYINPUT58), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n795_), .B2(new_n827_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n833_));
  OAI211_X1 g632(.A(new_n831_), .B(new_n758_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n823_), .A2(new_n826_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n538_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n823_), .A2(new_n826_), .A3(KEYINPUT119), .A4(new_n834_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n779_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n505_), .A2(new_n453_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n507_), .A2(new_n407_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT59), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n835_), .A2(new_n598_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n777_), .B(KEYINPUT54), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n848_));
  NAND2_X1  g647(.A1(new_n842_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n844_), .A2(new_n703_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G113gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n820_), .B2(new_n273_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n831_), .A2(new_n758_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n832_), .A2(new_n833_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n855_), .A2(new_n856_), .B1(new_n825_), .B2(new_n821_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n836_), .B1(new_n854_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n598_), .A3(new_n838_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n846_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n842_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n660_), .A2(G113gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n853_), .B1(new_n861_), .B2(new_n862_), .ZN(G1340gat));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n592_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n844_), .B2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n865_), .A2(KEYINPUT60), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT60), .ZN(new_n869_));
  AOI21_X1  g668(.A(G120gat), .B1(new_n659_), .B2(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n861_), .A2(new_n868_), .A3(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n864_), .B1(new_n867_), .B2(new_n871_), .ZN(new_n872_));
  OR4_X1    g671(.A1(new_n839_), .A2(new_n843_), .A3(new_n868_), .A4(new_n870_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n779_), .B1(new_n598_), .B2(new_n835_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n659_), .B1(new_n874_), .B2(new_n849_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n861_), .B2(KEYINPUT59), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n873_), .B(KEYINPUT121), .C1(new_n876_), .C2(new_n865_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n877_), .ZN(G1341gat));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n538_), .B2(KEYINPUT122), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(KEYINPUT122), .B2(new_n879_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n844_), .A2(new_n851_), .A3(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n861_), .B2(new_n598_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1342gat));
  NAND3_X1  g683(.A1(new_n844_), .A2(new_n758_), .A3(new_n851_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G134gat), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n273_), .A2(G134gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n861_), .B2(new_n887_), .ZN(G1343gat));
  NOR2_X1   g687(.A1(new_n839_), .A2(new_n635_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n624_), .A2(new_n408_), .A3(new_n453_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n561_), .A3(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT123), .B(G141gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1344gat));
  NAND3_X1  g692(.A1(new_n889_), .A2(new_n659_), .A3(new_n890_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT124), .B(G148gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1345gat));
  NAND2_X1  g695(.A1(new_n889_), .A2(new_n890_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n897_), .A2(new_n598_), .A3(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(new_n598_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1346gat));
  NAND4_X1  g700(.A1(new_n860_), .A2(new_n274_), .A3(new_n503_), .A4(new_n890_), .ZN(new_n902_));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT125), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n906_), .A3(new_n903_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n897_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n655_), .A2(new_n903_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n905_), .A2(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n505_), .A2(new_n407_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n635_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n644_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n847_), .A2(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n295_), .B1(new_n914_), .B2(new_n561_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n915_), .A2(KEYINPUT62), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n277_), .A3(new_n561_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(KEYINPUT62), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(G1348gat));
  NAND2_X1  g718(.A1(new_n914_), .A2(new_n659_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n839_), .A2(new_n454_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n912_), .A2(new_n296_), .A3(new_n592_), .ZN(new_n922_));
  AOI22_X1  g721(.A1(new_n920_), .A2(new_n276_), .B1(new_n921_), .B2(new_n922_), .ZN(G1349gat));
  NAND2_X1  g722(.A1(new_n847_), .A2(new_n913_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n924_), .A2(new_n292_), .A3(new_n598_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n921_), .A2(new_n635_), .A3(new_n538_), .A4(new_n911_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n281_), .ZN(G1350gat));
  NAND3_X1  g726(.A1(new_n914_), .A2(new_n274_), .A3(new_n293_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G190gat), .B1(new_n924_), .B2(new_n655_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT126), .ZN(G1351gat));
  NAND2_X1  g730(.A1(new_n911_), .A2(new_n454_), .ZN(new_n932_));
  AOI211_X1 g731(.A(new_n635_), .B(new_n932_), .C1(new_n859_), .C2(new_n846_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n561_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n659_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g736(.A(KEYINPUT63), .B(G211gat), .Z(new_n938_));
  AND3_X1   g737(.A1(new_n933_), .A2(new_n538_), .A3(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n933_), .A2(new_n538_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(G1354gat));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n943_), .B1(new_n933_), .B2(new_n758_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n932_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n273_), .A2(G218gat), .ZN(new_n946_));
  AND4_X1   g745(.A1(new_n503_), .A2(new_n860_), .A3(new_n945_), .A4(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(KEYINPUT127), .B1(new_n944_), .B2(new_n947_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n860_), .A2(new_n503_), .A3(new_n758_), .A4(new_n945_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(G218gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n933_), .A2(new_n946_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n948_), .A2(new_n953_), .ZN(G1355gat));
endmodule


