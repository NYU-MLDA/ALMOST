//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n971_, new_n972_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(KEYINPUT84), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(new_n208_), .B2(KEYINPUT84), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT85), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT84), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT85), .B1(new_n213_), .B2(new_n205_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(KEYINPUT87), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT3), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT2), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(new_n217_), .B2(new_n216_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n219_), .B(new_n221_), .C1(new_n218_), .C2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n217_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n220_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n225_), .A2(KEYINPUT1), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n227_), .B1(KEYINPUT1), .B2(new_n225_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n215_), .A2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n208_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n239_), .A2(KEYINPUT96), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(KEYINPUT96), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G1gat), .B(G29gat), .ZN(new_n245_));
  INV_X1    g044(.A(G85gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT4), .B1(new_n215_), .B2(new_n236_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(KEYINPUT4), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n243_), .B(KEYINPUT97), .Z(new_n254_));
  OAI211_X1 g053(.A(new_n244_), .B(new_n250_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT33), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n215_), .A2(new_n236_), .B1(KEYINPUT96), .B2(new_n239_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(new_n240_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n257_), .B1(new_n260_), .B2(new_n251_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT33), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n244_), .A4(new_n250_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n256_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n250_), .B1(new_n242_), .B2(new_n257_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n243_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(new_n253_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268_));
  INV_X1    g067(.A(G92gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT18), .B(G64gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n270_), .B(new_n271_), .Z(new_n272_));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT82), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(KEYINPUT24), .A3(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT25), .B(G183gat), .ZN(new_n277_));
  INV_X1    g076(.A(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT26), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(KEYINPUT26), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT95), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT23), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n274_), .B2(KEYINPUT24), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n276_), .A2(KEYINPUT95), .A3(new_n281_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n289_), .B1(KEYINPUT91), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT21), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(KEYINPUT21), .B2(new_n291_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n284_), .B1(G183gat), .B2(G190gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT22), .B(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n300_), .A3(new_n275_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n288_), .A2(new_n296_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n280_), .B(KEYINPUT81), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n277_), .A2(new_n279_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n276_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT83), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n285_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n276_), .B(KEYINPUT83), .C1(new_n304_), .C2(new_n305_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n303_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n302_), .B(KEYINPUT20), .C1(new_n310_), .C2(new_n296_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT19), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n288_), .A2(new_n301_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(new_n295_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n310_), .A2(new_n296_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n315_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n272_), .B1(new_n314_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n319_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n303_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT20), .B1(new_n323_), .B2(new_n296_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n313_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n272_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n325_), .B(new_n326_), .C1(new_n313_), .C2(new_n311_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n267_), .A2(new_n321_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n264_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n244_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n249_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n255_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n311_), .A2(new_n313_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n318_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n314_), .A2(new_n320_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n329_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT98), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n238_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n343_), .A2(KEYINPUT28), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(KEYINPUT28), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G22gat), .B(G50gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT90), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(new_n295_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT93), .ZN(new_n359_));
  XOR2_X1   g158(.A(G78gat), .B(G106gat), .Z(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n356_), .A3(new_n295_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT92), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n357_), .A2(KEYINPUT92), .A3(new_n356_), .A4(new_n295_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n360_), .B1(new_n359_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n354_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n360_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT93), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n358_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n365_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT94), .B1(new_n374_), .B2(new_n366_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n349_), .A2(new_n350_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT94), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n368_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n369_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n340_), .A2(new_n341_), .A3(new_n381_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n264_), .A2(new_n328_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT98), .B1(new_n383_), .B2(new_n380_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n374_), .A2(new_n366_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n378_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n376_), .B1(new_n374_), .B2(KEYINPUT94), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n332_), .B1(new_n388_), .B2(new_n369_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT99), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n308_), .A2(new_n309_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n301_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n316_), .B1(new_n392_), .B2(new_n295_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n315_), .B1(new_n393_), .B2(new_n302_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n322_), .A2(new_n324_), .A3(new_n313_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n272_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n390_), .B1(new_n396_), .B2(new_n327_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n334_), .A2(new_n335_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT99), .B1(new_n398_), .B2(new_n272_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT27), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n321_), .A2(new_n327_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n389_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n382_), .A2(new_n384_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G15gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(G71gat), .B(G99gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT30), .B(G43gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT86), .B1(new_n310_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n310_), .B2(new_n411_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n215_), .B(KEYINPUT31), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n414_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n332_), .ZN(new_n420_));
  AND4_X1   g219(.A1(new_n417_), .A2(new_n403_), .A3(new_n381_), .A4(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G15gat), .B(G22gat), .Z(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT75), .B(G8gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G1gat), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n426_), .B2(KEYINPUT14), .ZN(new_n427_));
  OR2_X1    g226(.A1(G1gat), .A2(G8gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G1gat), .A2(G8gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT76), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT76), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n432_), .A3(new_n429_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n427_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n433_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(new_n425_), .B2(G1gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n437_), .B2(new_n424_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G231gat), .A2(G233gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT11), .ZN(new_n442_));
  INV_X1    g241(.A(G57gat), .ZN(new_n443_));
  INV_X1    g242(.A(G64gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G57gat), .A2(G64gat), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT68), .ZN(new_n450_));
  AND2_X1   g249(.A1(G71gat), .A2(G78gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G71gat), .A2(G78gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n449_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n450_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n448_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(G57gat), .A2(G64gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G57gat), .A2(G64gat), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT11), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G71gat), .B(G78gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT68), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n449_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n447_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n456_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n441_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G127gat), .B(G155gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G183gat), .B(G211gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n465_), .A2(KEYINPUT17), .A3(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n470_), .B(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n454_), .A2(new_n455_), .A3(new_n448_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n447_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n456_), .A2(KEYINPUT69), .A3(new_n463_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n474_), .B1(new_n481_), .B2(new_n441_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(new_n441_), .B2(new_n481_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n472_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(G106gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT67), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n489_), .A2(KEYINPUT67), .A3(new_n490_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n493_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT66), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n269_), .A2(G85gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n246_), .A2(G92gat), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G85gat), .B(G92gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n502_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n485_), .B1(new_n501_), .B2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n489_), .A2(new_n496_), .A3(new_n497_), .A4(new_n490_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n503_), .A2(new_n504_), .A3(new_n502_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n511_), .B(new_n485_), .C1(new_n512_), .C2(new_n505_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT9), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G85gat), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n517_), .A2(new_n519_), .B1(new_n507_), .B2(new_n518_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT10), .B(G99gat), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n496_), .B(new_n497_), .C1(new_n521_), .C2(G106gat), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n520_), .A2(new_n522_), .A3(KEYINPUT65), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT65), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n519_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n518_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n487_), .A2(KEYINPUT10), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT10), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(G99gat), .ZN(new_n530_));
  AOI21_X1  g329(.A(G106gat), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(new_n498_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n524_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n533_));
  OAI22_X1  g332(.A1(new_n510_), .A2(new_n514_), .B1(new_n523_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535_));
  INV_X1    g334(.A(G29gat), .ZN(new_n536_));
  INV_X1    g335(.A(G36gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G29gat), .A2(G36gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G50gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(G50gat), .A3(new_n539_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT71), .B(G43gat), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n535_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n543_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n544_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(KEYINPUT15), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n534_), .A2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n498_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n555_), .A2(new_n500_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n513_), .B1(new_n556_), .B2(new_n485_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT65), .B1(new_n520_), .B2(new_n522_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n527_), .A2(new_n524_), .A3(new_n532_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n545_), .A2(new_n546_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT34), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT35), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n554_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n565_), .A2(new_n566_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G190gat), .B(G218gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT36), .ZN(new_n576_));
  INV_X1    g375(.A(new_n569_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n554_), .A2(new_n577_), .A3(new_n562_), .A4(new_n567_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n570_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n570_), .A2(KEYINPUT74), .A3(new_n576_), .A4(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n570_), .A2(new_n578_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n575_), .B(KEYINPUT36), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n484_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G120gat), .B(G148gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(G204gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT5), .B(G176gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n478_), .A2(new_n557_), .A3(new_n560_), .A4(new_n479_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n476_), .A2(new_n477_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n534_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT12), .B1(new_n480_), .B2(new_n534_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n479_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT69), .B1(new_n456_), .B2(new_n463_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n534_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n609_), .B2(new_n598_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n597_), .B1(new_n606_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n598_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n479_), .A2(new_n478_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n605_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n598_), .B(new_n601_), .C1(new_n613_), .C2(KEYINPUT12), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n614_), .B(new_n596_), .C1(new_n615_), .C2(new_n605_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n611_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT13), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(KEYINPUT70), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(KEYINPUT70), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n617_), .A2(new_n619_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n434_), .A2(new_n438_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n550_), .A2(KEYINPUT79), .A3(new_n551_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n630_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n547_), .A2(new_n552_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n634_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n631_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n439_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n630_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n629_), .B1(new_n638_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n641_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n637_), .B1(new_n644_), .B2(new_n634_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n553_), .A2(new_n630_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n646_), .A3(new_n636_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n629_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n643_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT80), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n626_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n420_), .A2(G1gat), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n423_), .A2(new_n592_), .A3(new_n652_), .A4(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT100), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n654_), .A2(new_n658_), .A3(new_n655_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n650_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n626_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n484_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n583_), .A2(new_n586_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n423_), .A2(new_n332_), .A3(new_n662_), .A4(new_n666_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(KEYINPUT101), .A3(G1gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT101), .B1(new_n667_), .B2(G1gat), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n659_), .A2(new_n660_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n202_), .B1(new_n657_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n656_), .B(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n659_), .A2(new_n660_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n668_), .A2(new_n669_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n673_), .A2(KEYINPUT103), .A3(new_n674_), .A4(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(G1324gat));
  AOI21_X1  g476(.A(new_n421_), .B1(new_n405_), .B2(new_n418_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n678_), .A2(new_n626_), .A3(new_n651_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n592_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n680_), .A2(new_n425_), .A3(new_n403_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n403_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n423_), .A2(new_n682_), .A3(new_n662_), .A4(new_n666_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  INV_X1    g485(.A(G8gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n685_), .A2(new_n686_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n686_), .B1(new_n685_), .B2(new_n688_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n681_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT40), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(KEYINPUT40), .B(new_n681_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1325gat));
  NAND2_X1  g494(.A1(new_n423_), .A2(new_n666_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n696_), .A2(new_n626_), .A3(new_n661_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n417_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G15gat), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(KEYINPUT41), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(KEYINPUT41), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n680_), .A2(G15gat), .A3(new_n418_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(G1326gat));
  INV_X1    g502(.A(G22gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n697_), .B2(new_n380_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT42), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n380_), .A2(new_n704_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n680_), .B2(new_n707_), .ZN(G1327gat));
  NOR2_X1   g507(.A1(new_n484_), .A2(new_n664_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n679_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n536_), .A3(new_n332_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n590_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n588_), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n678_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  INV_X1    g514(.A(new_n713_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n380_), .B1(new_n329_), .B2(new_n339_), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n717_), .A2(new_n341_), .B1(new_n389_), .B2(new_n403_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n417_), .B1(new_n718_), .B2(new_n384_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n715_), .B(new_n716_), .C1(new_n719_), .C2(new_n421_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n714_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n662_), .A2(new_n663_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT44), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n725_), .B(new_n722_), .C1(new_n714_), .C2(new_n720_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n724_), .A2(new_n726_), .A3(new_n420_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n711_), .B1(new_n727_), .B2(new_n536_), .ZN(G1328gat));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n724_), .A2(new_n726_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n537_), .B1(new_n730_), .B2(new_n682_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n679_), .A2(new_n537_), .A3(new_n682_), .A4(new_n709_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT45), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n731_), .B2(new_n734_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n724_), .A2(new_n726_), .A3(new_n403_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT46), .B(new_n733_), .C1(new_n736_), .C2(new_n537_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1329gat));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739_));
  INV_X1    g538(.A(G43gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n730_), .B2(new_n417_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n710_), .A2(new_n740_), .A3(new_n417_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n724_), .A2(new_n726_), .A3(new_n418_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT47), .B(new_n742_), .C1(new_n745_), .C2(new_n740_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1330gat));
  NAND2_X1  g546(.A1(new_n380_), .A2(new_n541_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT105), .Z(new_n749_));
  NAND2_X1  g548(.A1(new_n710_), .A2(new_n749_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n724_), .A2(new_n726_), .A3(new_n381_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n541_), .ZN(G1331gat));
  INV_X1    g551(.A(new_n626_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n678_), .A2(new_n753_), .A3(new_n650_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n592_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(KEYINPUT106), .A3(new_n592_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n332_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n651_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n696_), .A2(new_n753_), .A3(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n420_), .A2(new_n443_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n762_), .B2(new_n763_), .ZN(G1332gat));
  NAND4_X1  g563(.A1(new_n757_), .A2(new_n444_), .A3(new_n682_), .A4(new_n758_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT48), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n762_), .A2(new_n682_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G64gat), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT48), .B(new_n444_), .C1(new_n762_), .C2(new_n682_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT107), .B(new_n765_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1333gat));
  INV_X1    g573(.A(G71gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n762_), .B2(new_n417_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT49), .Z(new_n777_));
  NAND3_X1  g576(.A1(new_n759_), .A2(new_n775_), .A3(new_n417_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1334gat));
  INV_X1    g578(.A(G78gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n762_), .B2(new_n380_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT50), .Z(new_n782_));
  NAND3_X1  g581(.A1(new_n759_), .A2(new_n780_), .A3(new_n380_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1335gat));
  AND2_X1   g583(.A1(new_n754_), .A2(new_n709_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G85gat), .B1(new_n785_), .B2(new_n332_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n626_), .A2(new_n663_), .A3(new_n661_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT109), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n721_), .A2(KEYINPUT108), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n714_), .A2(new_n720_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n420_), .A2(new_n246_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n786_), .B1(new_n793_), .B2(new_n794_), .ZN(G1336gat));
  AOI21_X1  g594(.A(G92gat), .B1(new_n785_), .B2(new_n682_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n403_), .A2(new_n517_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n793_), .B2(new_n797_), .ZN(G1337gat));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799_));
  INV_X1    g598(.A(new_n521_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n785_), .A2(new_n800_), .A3(new_n417_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n793_), .A2(new_n417_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n799_), .B(new_n801_), .C1(new_n802_), .C2(new_n487_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n487_), .B1(new_n793_), .B2(new_n417_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n801_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT51), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(G1338gat));
  NAND3_X1  g606(.A1(new_n785_), .A2(new_n488_), .A3(new_n380_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n789_), .A2(new_n381_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n488_), .B1(new_n721_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n811_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n808_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT53), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n808_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1339gat));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n640_), .A2(new_n641_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n636_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n640_), .A2(new_n646_), .A3(new_n637_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n629_), .A3(new_n823_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n824_), .A2(new_n649_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n616_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n598_), .A2(new_n601_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n609_), .A2(new_n599_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n604_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n596_), .B1(new_n829_), .B2(new_n614_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n825_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n617_), .A2(KEYINPUT112), .A3(new_n825_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n604_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n829_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n827_), .A2(new_n828_), .A3(KEYINPUT55), .A4(new_n604_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(KEYINPUT56), .A4(new_n597_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n616_), .A2(new_n650_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n616_), .A2(new_n650_), .A3(KEYINPUT110), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n842_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n615_), .A2(new_n605_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n606_), .B1(KEYINPUT55), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n839_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n597_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n597_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(KEYINPUT111), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n835_), .B1(new_n848_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n820_), .B1(new_n857_), .B2(new_n665_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n820_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n842_), .A2(new_n847_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n597_), .ZN(new_n861_));
  AOI211_X1 g660(.A(new_n853_), .B(new_n596_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n863_), .B2(KEYINPUT111), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n664_), .B(new_n859_), .C1(new_n864_), .C2(new_n835_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n825_), .A2(new_n616_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n825_), .A2(KEYINPUT114), .A3(new_n616_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n713_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n870_), .B(KEYINPUT58), .C1(new_n862_), .C2(new_n861_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n858_), .A2(new_n865_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n663_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n878_));
  INV_X1    g677(.A(new_n625_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n761_), .B1(new_n879_), .B2(new_n623_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n592_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n651_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n591_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n877_), .A2(new_n884_), .ZN(new_n885_));
  NOR4_X1   g684(.A1(new_n682_), .A2(new_n418_), .A3(new_n380_), .A4(new_n420_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n885_), .A2(KEYINPUT115), .A3(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G113gat), .B1(new_n891_), .B2(new_n650_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n894_));
  MUX2_X1   g693(.A(new_n893_), .B(new_n894_), .S(new_n887_), .Z(new_n895_));
  AND2_X1   g694(.A1(new_n761_), .A2(G113gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n892_), .B1(new_n895_), .B2(new_n896_), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n753_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n891_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n895_), .A2(new_n626_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n898_), .ZN(G1341gat));
  XOR2_X1   g701(.A(KEYINPUT118), .B(G127gat), .Z(new_n903_));
  NAND3_X1  g702(.A1(new_n895_), .A2(new_n484_), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n663_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n907_));
  INV_X1    g706(.A(G127gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT117), .B1(new_n905_), .B2(G127gat), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n904_), .A2(new_n909_), .A3(new_n910_), .ZN(G1342gat));
  AOI21_X1  g710(.A(G134gat), .B1(new_n891_), .B2(new_n665_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n716_), .A2(G134gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT119), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n895_), .B2(new_n914_), .ZN(G1343gat));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n380_), .A2(new_n418_), .A3(new_n332_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n682_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n848_), .A2(new_n856_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n835_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n665_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n921_), .A2(new_n859_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n484_), .B1(new_n922_), .B2(new_n858_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n884_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n916_), .B(new_n918_), .C1(new_n923_), .C2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n876_), .B2(new_n663_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n918_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT120), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n925_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n650_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n626_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g732(.A1(new_n929_), .A2(new_n484_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT61), .B(G155gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1346gat));
  AOI21_X1  g735(.A(new_n916_), .B1(new_n885_), .B2(new_n918_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n926_), .A2(KEYINPUT120), .A3(new_n927_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n665_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(G162gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n939_), .A2(KEYINPUT121), .A3(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n664_), .B1(new_n925_), .B2(new_n928_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(G162gat), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n929_), .A2(G162gat), .A3(new_n716_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n941_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n941_), .A2(new_n944_), .A3(KEYINPUT122), .A4(new_n945_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1347gat));
  NOR2_X1   g749(.A1(new_n926_), .A2(new_n403_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n380_), .A2(new_n418_), .A3(new_n332_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n954_), .A2(new_n298_), .A3(new_n650_), .ZN(new_n955_));
  OAI21_X1  g754(.A(G169gat), .B1(new_n953_), .B2(new_n661_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n956_), .A2(new_n957_), .A3(KEYINPUT62), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n958_), .B1(new_n956_), .B2(KEYINPUT62), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n957_), .B1(new_n956_), .B2(KEYINPUT62), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n955_), .B1(new_n959_), .B2(new_n960_), .ZN(G1348gat));
  NOR2_X1   g760(.A1(new_n299_), .A2(KEYINPUT124), .ZN(new_n962_));
  XNOR2_X1  g761(.A(KEYINPUT124), .B(G176gat), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n953_), .A2(new_n753_), .ZN(new_n964_));
  MUX2_X1   g763(.A(new_n962_), .B(new_n963_), .S(new_n964_), .Z(G1349gat));
  NAND3_X1  g764(.A1(new_n954_), .A2(new_n484_), .A3(new_n277_), .ZN(new_n966_));
  OAI21_X1  g765(.A(G183gat), .B1(new_n953_), .B2(new_n663_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n968_), .B(new_n969_), .ZN(G1350gat));
  OAI21_X1  g769(.A(G190gat), .B1(new_n953_), .B2(new_n713_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n665_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n953_), .B2(new_n972_), .ZN(G1351gat));
  AND3_X1   g772(.A1(new_n951_), .A2(new_n418_), .A3(new_n389_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(new_n650_), .ZN(new_n975_));
  INV_X1    g774(.A(G197gat), .ZN(new_n976_));
  OR3_X1    g775(.A1(new_n975_), .A2(KEYINPUT126), .A3(new_n976_), .ZN(new_n977_));
  OAI21_X1  g776(.A(KEYINPUT126), .B1(new_n975_), .B2(new_n976_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n975_), .A2(new_n976_), .ZN(new_n979_));
  AND3_X1   g778(.A1(new_n977_), .A2(new_n978_), .A3(new_n979_), .ZN(G1352gat));
  NAND2_X1  g779(.A1(new_n974_), .A2(new_n626_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g781(.A1(new_n974_), .A2(new_n484_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(KEYINPUT63), .B(G211gat), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  INV_X1    g784(.A(KEYINPUT63), .ZN(new_n986_));
  INV_X1    g785(.A(G211gat), .ZN(new_n987_));
  NAND3_X1  g786(.A1(new_n983_), .A2(new_n986_), .A3(new_n987_), .ZN(new_n988_));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n988_), .A2(new_n989_), .ZN(new_n990_));
  NAND4_X1  g789(.A1(new_n983_), .A2(KEYINPUT127), .A3(new_n986_), .A4(new_n987_), .ZN(new_n991_));
  AOI21_X1  g790(.A(new_n985_), .B1(new_n990_), .B2(new_n991_), .ZN(G1354gat));
  AOI21_X1  g791(.A(G218gat), .B1(new_n974_), .B2(new_n665_), .ZN(new_n993_));
  AND2_X1   g792(.A1(new_n716_), .A2(G218gat), .ZN(new_n994_));
  AOI21_X1  g793(.A(new_n993_), .B1(new_n974_), .B2(new_n994_), .ZN(G1355gat));
endmodule


