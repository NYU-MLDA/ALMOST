//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(G204gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  OAI211_X1 g005(.A(KEYINPUT21), .B(new_n204_), .C1(new_n206_), .C2(new_n202_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G211gat), .B(G218gat), .Z(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n205_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT21), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT88), .ZN(new_n216_));
  NOR3_X1   g015(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT86), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT3), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT2), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n218_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n216_), .B1(new_n224_), .B2(KEYINPUT87), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT87), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n218_), .A2(new_n226_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(KEYINPUT1), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT84), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(KEYINPUT84), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT85), .ZN(new_n234_));
  OR3_X1    g033(.A1(new_n229_), .A2(new_n234_), .A3(KEYINPUT1), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(new_n229_), .B2(KEYINPUT1), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n220_), .A2(new_n222_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n228_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n214_), .B1(new_n240_), .B2(KEYINPUT29), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G22gat), .B(G50gat), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n225_), .A2(new_n227_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT28), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT29), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n247_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n245_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G78gat), .B(G106gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n246_), .A2(new_n248_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT28), .ZN(new_n256_));
  INV_X1    g055(.A(new_n245_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n249_), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n252_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n254_), .A2(KEYINPUT91), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n252_), .B2(new_n258_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n244_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n250_), .A2(new_n251_), .A3(new_n245_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n257_), .B1(new_n256_), .B2(new_n249_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n243_), .B(new_n259_), .C1(new_n266_), .C2(new_n261_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G169gat), .ZN(new_n270_));
  INV_X1    g069(.A(G176gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT81), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(G169gat), .B2(G176gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT82), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT24), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT25), .B(G183gat), .Z(new_n283_));
  INV_X1    g082(.A(G190gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT26), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(KEYINPUT80), .B2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G190gat), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT80), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT24), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n279_), .B(new_n289_), .C1(new_n277_), .C2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT22), .B(G169gat), .Z(new_n293_));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  OAI221_X1 g093(.A(new_n290_), .B1(new_n293_), .B2(G176gat), .C1(new_n282_), .C2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n214_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n277_), .A2(new_n291_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n282_), .B1(new_n278_), .B2(new_n275_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT92), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n287_), .B(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n301_), .B2(new_n283_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n295_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(new_n213_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT19), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n297_), .A2(KEYINPUT20), .A3(new_n304_), .A4(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n303_), .B2(new_n213_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n292_), .A2(new_n214_), .A3(new_n295_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n306_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G8gat), .B(G36gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n308_), .A2(new_n313_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT97), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT20), .B1(new_n303_), .B2(new_n213_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n306_), .B1(new_n322_), .B2(new_n296_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n312_), .B2(new_n306_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n318_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT97), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n308_), .A2(new_n313_), .A3(new_n326_), .A4(new_n319_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n321_), .A2(KEYINPUT27), .A3(new_n325_), .A4(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n322_), .A2(new_n296_), .A3(new_n306_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n307_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n318_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n320_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n328_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n269_), .A2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G1gat), .B(G29gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT94), .B(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT0), .B(G57gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G113gat), .B(G120gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n240_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n246_), .A2(new_n345_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT95), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n349_), .A2(KEYINPUT95), .A3(new_n350_), .A4(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n228_), .A2(new_n345_), .A3(new_n239_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n347_), .B1(new_n228_), .B2(new_n239_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT4), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n349_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n350_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n342_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n350_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n360_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n358_), .A2(KEYINPUT4), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n342_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n292_), .A2(new_n295_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT30), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n371_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(new_n347_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378_));
  INV_X1    g177(.A(G43gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT31), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n377_), .B(new_n381_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n337_), .A2(new_n370_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n369_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n349_), .A2(new_n364_), .A3(new_n351_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n342_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n359_), .A2(new_n361_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n350_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n332_), .A2(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n354_), .A2(new_n355_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n391_), .A2(KEYINPUT33), .A3(new_n368_), .A4(new_n367_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n329_), .A2(new_n330_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n324_), .B2(new_n395_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n370_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n269_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n268_), .B1(new_n393_), .B2(new_n398_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT96), .ZN(new_n404_));
  INV_X1    g203(.A(new_n370_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n336_), .A2(new_n405_), .A3(new_n268_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n383_), .B1(new_n407_), .B2(new_n382_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT74), .B(G1gat), .ZN(new_n409_));
  INV_X1    g208(.A(G8gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT14), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G15gat), .B(G22gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G1gat), .B(G8gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G29gat), .B(G36gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT72), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G43gat), .B(G50gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n419_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n418_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G229gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n422_), .A2(new_n426_), .A3(KEYINPUT15), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT15), .B1(new_n422_), .B2(new_n426_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n418_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n418_), .A2(new_n427_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n430_), .B1(new_n436_), .B2(new_n428_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G113gat), .B(G141gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT77), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G169gat), .B(G197gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(KEYINPUT78), .Z(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n444_), .B2(KEYINPUT79), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT79), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n446_), .B(new_n443_), .C1(new_n435_), .C2(new_n437_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n408_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(KEYINPUT71), .ZN(new_n451_));
  AND2_X1   g250(.A1(G230gat), .A2(G233gat), .ZN(new_n452_));
  OR2_X1    g251(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n453_));
  INV_X1    g252(.A(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT64), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT64), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n453_), .A2(new_n455_), .A3(new_n457_), .A4(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(KEYINPUT9), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G85gat), .ZN(new_n466_));
  INV_X1    g265(.A(G92gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT9), .A3(new_n463_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n459_), .A2(new_n462_), .A3(new_n465_), .A4(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT65), .ZN(new_n471_));
  AND2_X1   g270(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT64), .B(G106gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n464_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n462_), .A4(new_n469_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n471_), .A2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT66), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n485_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n488_));
  INV_X1    g287(.A(G99gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n454_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(KEYINPUT8), .B(new_n482_), .C1(new_n487_), .C2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n482_), .B1(new_n487_), .B2(new_n495_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n479_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(KEYINPUT11), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n505_));
  XOR2_X1   g304(.A(G71gat), .B(G78gat), .Z(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(KEYINPUT11), .B2(new_n502_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n507_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n509_), .B1(new_n510_), .B2(new_n503_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n452_), .B1(new_n500_), .B2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n470_), .A2(KEYINPUT65), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT9), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n480_), .A2(new_n481_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n493_), .A2(new_n494_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n477_), .B1(new_n518_), .B2(new_n476_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n496_), .B(new_n499_), .C1(new_n514_), .C2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n508_), .A2(new_n511_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n508_), .A2(new_n511_), .A3(KEYINPUT68), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT68), .B1(new_n508_), .B2(new_n511_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n520_), .B(KEYINPUT12), .C1(new_n525_), .C2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n513_), .A2(new_n524_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n522_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n520_), .A2(new_n521_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n452_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT69), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n528_), .A2(new_n531_), .A3(KEYINPUT69), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G120gat), .B(G148gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G176gat), .B(G204gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n528_), .A2(new_n531_), .A3(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(KEYINPUT70), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n534_), .A2(new_n544_), .A3(new_n535_), .A4(new_n539_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n451_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n450_), .A2(KEYINPUT71), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n418_), .B(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n525_), .A2(new_n526_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT76), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(new_n554_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n553_), .A2(new_n521_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n553_), .A2(new_n521_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n559_), .B(KEYINPUT17), .Z(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n520_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  OAI221_X1 g371(.A(new_n570_), .B1(KEYINPUT35), .B2(new_n572_), .C1(new_n520_), .C2(new_n427_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(KEYINPUT35), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT73), .ZN(new_n579_));
  XOR2_X1   g378(.A(G134gat), .B(G162gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n573_), .A2(new_n575_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n576_), .A2(new_n577_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n581_), .B(KEYINPUT36), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n584_), .A2(KEYINPUT37), .A3(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT37), .B1(new_n584_), .B2(new_n587_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n569_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n449_), .A2(new_n551_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n370_), .A3(new_n409_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT38), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT99), .B1(new_n584_), .B2(new_n587_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n587_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(new_n583_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n408_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n550_), .A2(new_n569_), .A3(new_n448_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n370_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n604_), .A2(KEYINPUT101), .A3(G1gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT101), .B1(new_n604_), .B2(G1gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n593_), .B1(new_n605_), .B2(new_n606_), .ZN(G1324gat));
  NAND3_X1  g406(.A1(new_n591_), .A2(new_n410_), .A3(new_n335_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n599_), .A2(new_n335_), .A3(new_n601_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n609_), .A2(new_n610_), .A3(G8gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n609_), .B2(G8gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(G1325gat));
  NOR2_X1   g414(.A1(new_n602_), .A2(new_n603_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G15gat), .B1(new_n616_), .B2(new_n382_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(KEYINPUT41), .ZN(new_n618_));
  INV_X1    g417(.A(new_n382_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n591_), .A2(new_n373_), .A3(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT103), .Z(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(KEYINPUT41), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n618_), .A2(new_n621_), .A3(new_n622_), .ZN(G1326gat));
  INV_X1    g422(.A(G22gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n591_), .A2(new_n624_), .A3(new_n268_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n268_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n626_));
  XOR2_X1   g425(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n627_));
  AND3_X1   g426(.A1(new_n626_), .A2(G22gat), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n626_), .B2(G22gat), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n625_), .B1(new_n628_), .B2(new_n629_), .ZN(G1327gat));
  INV_X1    g429(.A(new_n598_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n569_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n550_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n449_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G29gat), .B1(new_n635_), .B2(new_n370_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n550_), .A2(new_n632_), .A3(new_n448_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n406_), .B1(new_n403_), .B2(KEYINPUT96), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n401_), .B(new_n268_), .C1(new_n398_), .C2(new_n393_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n382_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n383_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n588_), .A2(new_n589_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n638_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT43), .B(new_n644_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n637_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT44), .B(new_n637_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n370_), .A2(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n636_), .B1(new_n652_), .B2(new_n653_), .ZN(G1328gat));
  XNOR2_X1  g453(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(new_n651_), .A3(new_n335_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G36gat), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n336_), .A2(G36gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n635_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT45), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n656_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n661_), .B(KEYINPUT45), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n658_), .A3(new_n655_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1329gat));
  NOR2_X1   g466(.A1(new_n382_), .A2(new_n379_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n650_), .A2(new_n651_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT106), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n650_), .A2(new_n651_), .A3(new_n671_), .A4(new_n668_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n379_), .B1(new_n634_), .B2(new_n382_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n670_), .A2(new_n672_), .A3(new_n673_), .A4(new_n675_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1330gat));
  AOI21_X1  g478(.A(G50gat), .B1(new_n635_), .B2(new_n268_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n268_), .A2(G50gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n652_), .B2(new_n681_), .ZN(G1331gat));
  INV_X1    g481(.A(new_n448_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n569_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n599_), .A2(new_n550_), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n405_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n408_), .A2(new_n683_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n550_), .A3(new_n590_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT108), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n405_), .A2(G57gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(G1332gat));
  OAI21_X1  g490(.A(G64gat), .B1(new_n685_), .B2(new_n336_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT48), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT48), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n336_), .A2(G64gat), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n693_), .A2(new_n694_), .B1(new_n689_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI221_X1 g497(.A(KEYINPUT109), .B1(new_n689_), .B2(new_n695_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1333gat));
  OR2_X1    g499(.A1(new_n685_), .A2(new_n382_), .ZN(new_n701_));
  XOR2_X1   g500(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(G71gat), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(G71gat), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n382_), .A2(G71gat), .ZN(new_n705_));
  OAI22_X1  g504(.A1(new_n703_), .A2(new_n704_), .B1(new_n689_), .B2(new_n705_), .ZN(G1334gat));
  OAI21_X1  g505(.A(G78gat), .B1(new_n685_), .B2(new_n269_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT50), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n269_), .A2(G78gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n689_), .B2(new_n709_), .ZN(G1335gat));
  NOR2_X1   g509(.A1(new_n631_), .A2(new_n632_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n687_), .A2(new_n550_), .A3(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(new_n466_), .A3(new_n370_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n550_), .A2(new_n569_), .A3(new_n448_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n408_), .B2(new_n644_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n643_), .A2(new_n638_), .A3(new_n645_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT111), .Z(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n370_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n713_), .B1(new_n719_), .B2(new_n466_), .ZN(G1336gat));
  AOI21_X1  g519(.A(G92gat), .B1(new_n712_), .B2(new_n335_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT112), .Z(new_n722_));
  NOR2_X1   g521(.A1(new_n336_), .A2(new_n467_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n718_), .B2(new_n723_), .ZN(G1337gat));
  NOR3_X1   g523(.A1(new_n382_), .A2(new_n473_), .A3(new_n472_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n687_), .A2(new_n550_), .A3(new_n711_), .A4(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT113), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n489_), .B1(new_n717_), .B2(new_n619_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(G1338gat));
  NAND2_X1  g530(.A1(new_n717_), .A2(new_n268_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G106gat), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n268_), .A2(new_n475_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n687_), .A2(new_n550_), .A3(new_n711_), .A4(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT115), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n736_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT53), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n735_), .A2(new_n742_), .A3(new_n736_), .A4(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1339gat));
  NAND4_X1  g543(.A1(new_n590_), .A2(new_n549_), .A3(new_n548_), .A4(new_n448_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT54), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT117), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n435_), .A2(new_n437_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n436_), .A2(new_n428_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n441_), .B1(new_n749_), .B2(new_n429_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n434_), .B(new_n430_), .C1(new_n427_), .C2(new_n418_), .ZN(new_n751_));
  AOI22_X1  g550(.A1(new_n748_), .A2(new_n441_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n528_), .A2(KEYINPUT69), .A3(new_n531_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT69), .B1(new_n528_), .B2(new_n531_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n541_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n542_), .A2(KEYINPUT70), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n545_), .B(new_n752_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT116), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n543_), .A2(new_n759_), .A3(new_n545_), .A4(new_n752_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n542_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n524_), .A2(new_n527_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n452_), .B1(new_n763_), .B2(new_n530_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n528_), .A2(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n513_), .A2(new_n524_), .A3(new_n527_), .A4(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n539_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT56), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n539_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n762_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n761_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n594_), .A2(KEYINPUT57), .A3(new_n597_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n747_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n773_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n779_), .A2(new_n776_), .A3(KEYINPUT117), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n771_), .A2(new_n772_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n752_), .A2(new_n542_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n782_), .A2(KEYINPUT58), .A3(new_n783_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n645_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n779_), .B2(new_n598_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n781_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n746_), .B1(new_n792_), .B2(new_n632_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n619_), .A2(new_n370_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(new_n337_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n793_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n781_), .B2(new_n791_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n775_), .A2(new_n747_), .A3(new_n777_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT117), .B1(new_n779_), .B2(new_n776_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n803_), .A2(KEYINPUT118), .A3(new_n790_), .A4(new_n788_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n569_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n796_), .B1(new_n805_), .B2(new_n746_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n683_), .B(new_n798_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(G113gat), .ZN(new_n809_));
  INV_X1    g608(.A(G113gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n810_), .A3(new_n683_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT119), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n809_), .A2(new_n814_), .A3(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(G1340gat));
  OAI211_X1 g615(.A(new_n550_), .B(new_n798_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G120gat), .ZN(new_n818_));
  INV_X1    g617(.A(G120gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n551_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n806_), .B(new_n820_), .C1(KEYINPUT60), .C2(new_n819_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n818_), .A2(KEYINPUT120), .A3(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n806_), .A2(new_n827_), .A3(new_n632_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n806_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n829_), .A2(KEYINPUT59), .B1(new_n793_), .B2(new_n797_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n632_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n832_), .B2(new_n827_), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n829_), .B2(new_n631_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n836_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n644_), .A2(new_n834_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n837_), .A2(new_n838_), .B1(new_n830_), .B2(new_n839_), .ZN(G1343gat));
  NAND2_X1  g639(.A1(new_n805_), .A2(new_n746_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n619_), .A2(new_n269_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n405_), .A2(new_n335_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n683_), .A3(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n550_), .A3(new_n844_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g647(.A1(new_n843_), .A2(new_n632_), .A3(new_n844_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1346gat));
  NAND2_X1  g650(.A1(new_n843_), .A2(new_n844_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G162gat), .B1(new_n852_), .B2(new_n644_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n631_), .A2(G162gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n852_), .B2(new_n854_), .ZN(G1347gat));
  NOR2_X1   g654(.A1(new_n336_), .A2(new_n370_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(new_n268_), .A3(new_n382_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n793_), .A2(new_n683_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(G169gat), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n859_), .A2(new_n293_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT122), .ZN(G1348gat));
  NAND2_X1  g665(.A1(new_n841_), .A2(new_n269_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n867_), .A2(KEYINPUT124), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n857_), .A2(new_n382_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(KEYINPUT124), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n551_), .A2(new_n271_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n793_), .A2(new_n858_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n271_), .B1(new_n873_), .B2(new_n551_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n874_), .A2(new_n875_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n871_), .A2(new_n872_), .B1(new_n876_), .B2(new_n877_), .ZN(G1349gat));
  INV_X1    g677(.A(new_n283_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n873_), .A2(new_n879_), .A3(new_n569_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT125), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n868_), .A2(new_n632_), .A3(new_n869_), .A4(new_n870_), .ZN(new_n882_));
  INV_X1    g681(.A(G183gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n873_), .B2(new_n644_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n631_), .A2(new_n301_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n873_), .B2(new_n886_), .ZN(G1351gat));
  AND3_X1   g686(.A1(new_n841_), .A2(new_n842_), .A3(new_n856_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n683_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n550_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n569_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n888_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT126), .Z(new_n897_));
  OAI21_X1  g696(.A(new_n893_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n897_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n888_), .A2(KEYINPUT127), .A3(new_n899_), .A4(new_n894_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n897_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n898_), .A2(new_n900_), .A3(new_n901_), .ZN(G1354gat));
  INV_X1    g701(.A(new_n888_), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n903_), .A2(G218gat), .A3(new_n631_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G218gat), .B1(new_n903_), .B2(new_n644_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1355gat));
endmodule


