//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n204_), .B1(G99gat), .B2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT10), .B(G99gat), .Z(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n212_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n214_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n219_), .B(new_n216_), .C1(new_n208_), .C2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT64), .B1(new_n205_), .B2(new_n207_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n222_), .A2(new_n223_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n226_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n219_), .B1(new_n232_), .B2(new_n216_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n225_), .B1(new_n233_), .B2(KEYINPUT65), .ZN(new_n234_));
  INV_X1    g033(.A(new_n216_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n229_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(new_n224_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n237_), .B2(new_n230_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n219_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n218_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G29gat), .B(G36gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n242_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT15), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT15), .ZN(new_n251_));
  INV_X1    g050(.A(new_n249_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(new_n247_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n241_), .A2(new_n250_), .A3(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n239_), .B1(new_n238_), .B2(new_n219_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n232_), .A2(new_n216_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n257_), .A3(new_n225_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n258_), .B(new_n218_), .C1(new_n252_), .C2(new_n247_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G232gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT34), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n254_), .B(new_n259_), .C1(KEYINPUT35), .C2(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n261_), .A2(KEYINPUT35), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n253_), .A2(new_n250_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n218_), .B2(new_n258_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n263_), .B1(new_n265_), .B2(KEYINPUT71), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n254_), .A2(new_n259_), .A3(KEYINPUT71), .A4(new_n263_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G190gat), .B(G218gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G134gat), .B(G162gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(KEYINPUT36), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n203_), .B1(new_n269_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n273_), .ZN(new_n275_));
  AOI211_X1 g074(.A(KEYINPUT72), .B(new_n275_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n272_), .B(KEYINPUT36), .Z(new_n278_));
  NAND3_X1  g077(.A1(new_n267_), .A2(new_n268_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT73), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n267_), .A2(new_n281_), .A3(new_n268_), .A4(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n202_), .B1(new_n277_), .B2(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(KEYINPUT37), .B(new_n279_), .C1(new_n274_), .C2(new_n276_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G15gat), .B(G22gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT74), .B(G1gat), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n289_), .A2(G8gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT14), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n288_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G8gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G231gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT75), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n294_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G57gat), .B(G64gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G71gat), .B(G78gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT11), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n298_), .A2(KEYINPUT11), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(new_n299_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n298_), .A2(KEYINPUT11), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n297_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G155gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT16), .ZN(new_n307_));
  XOR2_X1   g106(.A(G183gat), .B(G211gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n305_), .B1(KEYINPUT17), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n309_), .B(KEYINPUT17), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n313_), .B2(new_n305_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n287_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT76), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G230gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n304_), .B(new_n218_), .C1(new_n234_), .C2(new_n240_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n258_), .A2(KEYINPUT66), .A3(new_n304_), .A4(new_n218_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n304_), .B1(new_n258_), .B2(new_n218_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n319_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n320_), .A2(new_n318_), .ZN(new_n327_));
  AOI211_X1 g126(.A(KEYINPUT12), .B(new_n304_), .C1(new_n258_), .C2(new_n218_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT12), .ZN(new_n329_));
  INV_X1    g128(.A(new_n304_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n241_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n327_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G120gat), .B(G148gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(G176gat), .B(G204gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n326_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n337_), .B(KEYINPUT68), .Z(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n326_), .B2(new_n332_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT13), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(KEYINPUT13), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n252_), .B2(new_n247_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n248_), .A2(KEYINPUT77), .A3(new_n249_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n294_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n294_), .A2(new_n253_), .A3(new_n250_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G229gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT78), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n349_), .A2(new_n350_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n294_), .B1(new_n348_), .B2(new_n347_), .ZN(new_n359_));
  OAI211_X1 g158(.A(G229gat), .B(G233gat), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n351_), .A2(KEYINPUT79), .A3(new_n352_), .A4(new_n354_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G113gat), .B(G141gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G169gat), .B(G197gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(KEYINPUT80), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n357_), .A2(new_n360_), .A3(new_n368_), .A4(new_n361_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n345_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT20), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n373_));
  INV_X1    g172(.A(G169gat), .ZN(new_n374_));
  INV_X1    g173(.A(G176gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n376_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n373_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT26), .B(G190gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT25), .B(G183gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n384_), .A2(KEYINPUT93), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT93), .B1(new_n384_), .B2(new_n387_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n381_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT22), .B(G169gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n375_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n382_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n378_), .B(KEYINPUT23), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(G183gat), .B2(G190gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT94), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT94), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n399_), .A3(new_n396_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n390_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(G197gat), .A2(G204gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT21), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(KEYINPUT21), .A3(new_n403_), .ZN(new_n407_));
  INV_X1    g206(.A(G211gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT90), .B1(new_n408_), .B2(G218gat), .ZN(new_n409_));
  INV_X1    g208(.A(G218gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(G211gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n406_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G197gat), .B(G204gat), .Z(new_n414_));
  OAI211_X1 g213(.A(new_n414_), .B(KEYINPUT21), .C1(new_n411_), .C2(new_n409_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n372_), .B1(new_n401_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n395_), .B1(KEYINPUT24), .B2(new_n376_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(KEYINPUT24), .B2(new_n383_), .ZN(new_n419_));
  INV_X1    g218(.A(G183gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT25), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT83), .B(G190gat), .Z(new_n422_));
  INV_X1    g221(.A(KEYINPUT26), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n421_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n427_));
  NOR2_X1   g226(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n428_));
  OAI21_X1  g227(.A(G183gat), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT82), .Z(new_n430_));
  OAI21_X1  g229(.A(new_n419_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n394_), .A2(KEYINPUT84), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n422_), .A2(new_n420_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n395_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n393_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n431_), .A2(new_n415_), .A3(new_n437_), .A4(new_n413_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n417_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT19), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n431_), .A2(new_n437_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n416_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n441_), .A2(new_n372_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n444_), .B(new_n445_), .C1(new_n416_), .C2(new_n401_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT18), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT27), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT102), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n451_), .B(KEYINPUT101), .Z(new_n456_));
  INV_X1    g255(.A(KEYINPUT99), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n413_), .A2(KEYINPUT91), .A3(new_n415_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT91), .B1(new_n413_), .B2(new_n415_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n390_), .B(new_n397_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n444_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT98), .B1(new_n460_), .B2(KEYINPUT20), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n441_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n441_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n417_), .A2(new_n465_), .A3(new_n438_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n457_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n390_), .A2(new_n397_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n458_), .A2(new_n459_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT20), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT98), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n461_), .A3(new_n444_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT99), .B1(new_n474_), .B2(new_n441_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n455_), .B(new_n456_), .C1(new_n468_), .C2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n464_), .A2(new_n457_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n466_), .B1(new_n474_), .B2(new_n441_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n457_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n455_), .B1(new_n480_), .B2(new_n456_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n454_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G22gat), .B(G50gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G155gat), .A2(G162gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G155gat), .A2(G162gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G141gat), .A2(G148gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT3), .Z(new_n491_));
  NAND2_X1  g290(.A1(G141gat), .A2(G148gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT2), .Z(new_n493_));
  OAI211_X1 g292(.A(new_n487_), .B(new_n489_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n488_), .B1(KEYINPUT1), .B2(new_n487_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(KEYINPUT1), .B2(new_n487_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n490_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n492_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT29), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n470_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(G228gat), .A3(G233gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G228gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT89), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n416_), .B(new_n505_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n500_), .A2(new_n501_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT28), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n507_), .A2(new_n509_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n486_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n510_), .A3(new_n485_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n447_), .A2(new_n452_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n451_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(KEYINPUT27), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G225gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G127gat), .B(G134gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G113gat), .B(G120gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n525_), .B(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n500_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n499_), .A2(new_n532_), .A3(new_n530_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n524_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(KEYINPUT4), .A3(new_n535_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n533_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT4), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n538_), .A2(KEYINPUT95), .A3(new_n539_), .A4(new_n499_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT95), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n541_), .B1(new_n535_), .B2(KEYINPUT4), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n536_), .B1(new_n543_), .B2(new_n524_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G57gat), .B(G85gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT97), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(G1gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n548_));
  INV_X1    g347(.A(G29gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n547_), .B(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT100), .B1(new_n544_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n543_), .A2(new_n524_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n536_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n553_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n544_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n551_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n557_), .A2(KEYINPUT100), .A3(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G227gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT85), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT30), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G15gat), .B(G43gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G71gat), .B(G99gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n443_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n443_), .A2(new_n568_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n565_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n564_), .A3(new_n569_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n561_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n533_), .B(KEYINPUT31), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n572_), .A2(new_n574_), .A3(new_n561_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n576_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n580_), .B2(new_n575_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n560_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n482_), .A2(new_n517_), .A3(new_n522_), .A4(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT103), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n456_), .B1(new_n468_), .B2(new_n475_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT102), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n476_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n521_), .B1(new_n588_), .B2(new_n454_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n589_), .A2(KEYINPUT103), .A3(new_n517_), .A4(new_n582_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n453_), .B1(new_n587_), .B2(new_n476_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n516_), .B1(new_n559_), .B2(new_n556_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n592_), .A2(new_n593_), .A3(new_n521_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n451_), .A2(KEYINPUT32), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n480_), .A2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n560_), .B(new_n596_), .C1(new_n595_), .C2(new_n447_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n544_), .A2(new_n551_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n534_), .A2(new_n535_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n558_), .B1(new_n600_), .B2(new_n524_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n543_), .A2(new_n524_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n598_), .A2(KEYINPUT33), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n603_), .B(new_n520_), .C1(KEYINPUT33), .C2(new_n598_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n516_), .B1(new_n597_), .B2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n581_), .B1(new_n594_), .B2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n371_), .B1(new_n591_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n317_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n560_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n608_), .A2(new_n289_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n371_), .A2(new_n314_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT104), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n277_), .A2(new_n283_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n591_), .B2(new_n606_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(new_n609_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n610_), .A2(new_n611_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n612_), .A2(new_n619_), .A3(new_n620_), .ZN(G1324gat));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622_));
  INV_X1    g421(.A(new_n589_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G8gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT105), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n627_), .A3(G8gat), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n626_), .A2(KEYINPUT39), .A3(new_n628_), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n608_), .A2(G8gat), .A3(new_n589_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n626_), .B2(KEYINPUT39), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n622_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n626_), .A2(KEYINPUT39), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n626_), .A2(KEYINPUT39), .A3(new_n628_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n633_), .A2(KEYINPUT40), .A3(new_n634_), .A4(new_n630_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n581_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n617_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n637_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n608_), .B2(new_n641_), .ZN(G1326gat));
  OAI21_X1  g441(.A(G22gat), .B1(new_n618_), .B2(new_n517_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT42), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n517_), .A2(G22gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n608_), .B2(new_n645_), .ZN(G1327gat));
  NAND2_X1  g445(.A1(new_n615_), .A2(new_n314_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT107), .Z(new_n648_));
  AND2_X1   g447(.A1(new_n607_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n560_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n371_), .A2(new_n315_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT106), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n286_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n591_), .A2(new_n606_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(new_n286_), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n287_), .B(new_n654_), .C1(new_n591_), .C2(new_n606_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n651_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT44), .B(new_n651_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n609_), .A2(new_n549_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n650_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n649_), .A2(new_n666_), .A3(new_n623_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT45), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(new_n623_), .A3(new_n662_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(G36gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G36gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n668_), .B(new_n674_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1329gat));
  NAND3_X1  g477(.A1(new_n663_), .A2(G43gat), .A3(new_n638_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT110), .B(G43gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n649_), .B2(new_n638_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g483(.A(G50gat), .B1(new_n649_), .B2(new_n516_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n516_), .A2(G50gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n663_), .B2(new_n686_), .ZN(G1331gat));
  NOR2_X1   g486(.A1(new_n345_), .A2(new_n370_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n616_), .A2(new_n315_), .A3(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G57gat), .B1(new_n689_), .B2(new_n609_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n656_), .A2(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n317_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n609_), .A2(G57gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(G1332gat));
  OAI21_X1  g493(.A(G64gat), .B1(new_n689_), .B2(new_n589_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT48), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n589_), .A2(G64gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n692_), .B2(new_n697_), .ZN(G1333gat));
  OAI21_X1  g497(.A(G71gat), .B1(new_n689_), .B2(new_n581_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT49), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n581_), .A2(G71gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n692_), .B2(new_n701_), .ZN(G1334gat));
  OAI21_X1  g501(.A(G78gat), .B1(new_n689_), .B2(new_n517_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT50), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n517_), .A2(G78gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n692_), .B2(new_n705_), .ZN(G1335gat));
  NAND2_X1  g505(.A1(new_n691_), .A2(new_n648_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n209_), .B1(new_n707_), .B2(new_n609_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT111), .Z(new_n709_));
  OR2_X1    g508(.A1(new_n657_), .A2(new_n658_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n710_), .A2(new_n314_), .A3(new_n688_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n609_), .A2(new_n209_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1336gat));
  AND2_X1   g512(.A1(new_n711_), .A2(new_n623_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n623_), .A2(new_n210_), .ZN(new_n715_));
  OAI22_X1  g514(.A1(new_n714_), .A2(new_n210_), .B1(new_n707_), .B2(new_n715_), .ZN(G1337gat));
  AND4_X1   g515(.A1(new_n213_), .A2(new_n691_), .A3(new_n638_), .A4(new_n648_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n711_), .A2(new_n638_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n221_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT51), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n722_), .B(new_n718_), .C1(new_n719_), .C2(new_n221_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1338gat));
  NOR3_X1   g523(.A1(new_n707_), .A2(G106gat), .A3(new_n517_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT112), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n710_), .A2(new_n314_), .A3(new_n516_), .A4(new_n688_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G106gat), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n726_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n726_), .A2(new_n730_), .A3(new_n734_), .A4(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1339gat));
  INV_X1    g535(.A(KEYINPUT119), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n343_), .A2(new_n344_), .ZN(new_n738_));
  OR4_X1    g537(.A1(new_n314_), .A2(new_n286_), .A3(new_n370_), .A4(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n354_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n358_), .A2(new_n359_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n354_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  MUX2_X1   g544(.A(new_n745_), .B(new_n362_), .S(new_n365_), .Z(new_n746_));
  NOR2_X1   g545(.A1(new_n328_), .A2(new_n331_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n319_), .B1(new_n747_), .B2(new_n324_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n332_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n327_), .B(KEYINPUT55), .C1(new_n328_), .C2(new_n331_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n748_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n340_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(KEYINPUT56), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT56), .B1(new_n752_), .B2(new_n753_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n338_), .B(new_n746_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(KEYINPUT58), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n758_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n286_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n754_), .A2(new_n755_), .A3(KEYINPUT113), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n752_), .A2(new_n753_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(KEYINPUT113), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n370_), .A2(new_n338_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n763_), .B1(new_n764_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n765_), .A2(new_n766_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n752_), .A2(KEYINPUT56), .A3(new_n753_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n768_), .B1(new_n755_), .B2(KEYINPUT113), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(KEYINPUT114), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n746_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT115), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n746_), .B(new_n780_), .C1(new_n341_), .C2(new_n339_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n771_), .A2(new_n777_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n615_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(KEYINPUT57), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n762_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n784_), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n785_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n775_), .A2(new_n776_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n782_), .B1(new_n791_), .B2(new_n763_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n615_), .B1(new_n792_), .B2(new_n777_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n784_), .A2(new_n785_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT116), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n788_), .B(new_n789_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n741_), .B1(new_n798_), .B2(new_n314_), .ZN(new_n799_));
  NOR4_X1   g598(.A1(new_n623_), .A2(new_n609_), .A3(new_n516_), .A4(new_n581_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n737_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n786_), .A2(new_n787_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n803_), .A2(new_n789_), .A3(new_n761_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT57), .B1(new_n796_), .B2(KEYINPUT116), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(KEYINPUT116), .B2(new_n796_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n315_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT119), .B(new_n800_), .C1(new_n807_), .C2(new_n741_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n802_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(G113gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n370_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n795_), .A2(new_n797_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n803_), .A2(new_n789_), .A3(new_n761_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n314_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n741_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n816_), .B(new_n800_), .C1(KEYINPUT120), .C2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n370_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(G113gat), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n811_), .A2(new_n823_), .ZN(G1340gat));
  NAND3_X1  g623(.A1(new_n818_), .A2(new_n738_), .A3(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G120gat), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n345_), .A2(KEYINPUT60), .ZN(new_n827_));
  MUX2_X1   g626(.A(new_n827_), .B(KEYINPUT60), .S(G120gat), .Z(new_n828_));
  NAND2_X1  g627(.A1(new_n809_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(G1341gat));
  NAND2_X1  g629(.A1(new_n809_), .A2(new_n315_), .ZN(new_n831_));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n818_), .A2(new_n821_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n314_), .A2(new_n832_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT121), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n831_), .A2(new_n832_), .B1(new_n833_), .B2(new_n835_), .ZN(G1342gat));
  AND4_X1   g635(.A1(G134gat), .A2(new_n818_), .A3(new_n286_), .A4(new_n821_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n802_), .A2(new_n808_), .A3(new_n615_), .ZN(new_n838_));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT122), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n842_), .A3(new_n839_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n837_), .B1(new_n841_), .B2(new_n843_), .ZN(G1343gat));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845_));
  NOR4_X1   g644(.A1(new_n623_), .A2(new_n609_), .A3(new_n517_), .A4(new_n638_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n816_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n816_), .B2(new_n846_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n370_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g649(.A(new_n738_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g651(.A(new_n315_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1346gat));
  INV_X1    g654(.A(G162gat), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n615_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n847_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n848_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n287_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n857_), .B1(new_n860_), .B2(new_n856_), .ZN(G1347gat));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n623_), .A2(new_n370_), .A3(new_n582_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT124), .Z(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n799_), .A2(new_n516_), .A3(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n866_), .A2(KEYINPUT125), .A3(new_n374_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n816_), .A2(new_n517_), .A3(new_n864_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(G169gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n862_), .B1(new_n867_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n816_), .A2(new_n517_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n623_), .A2(new_n582_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n370_), .A3(new_n391_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT125), .B1(new_n866_), .B2(new_n374_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n869_), .A2(new_n868_), .A3(G169gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(KEYINPUT62), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n871_), .A2(new_n875_), .A3(new_n878_), .ZN(G1348gat));
  NAND2_X1  g678(.A1(new_n874_), .A2(new_n738_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g680(.A1(new_n420_), .A2(KEYINPUT126), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n874_), .A2(new_n315_), .A3(new_n386_), .A4(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n874_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n314_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(KEYINPUT126), .A2(G183gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n885_), .B2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n884_), .B2(new_n287_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n874_), .A2(new_n615_), .A3(new_n385_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1351gat));
  NAND3_X1  g689(.A1(new_n609_), .A2(new_n516_), .A3(new_n581_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n891_), .A2(KEYINPUT127), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(KEYINPUT127), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n799_), .A2(new_n589_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n370_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n738_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n315_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  NAND3_X1  g703(.A1(new_n895_), .A2(new_n410_), .A3(new_n615_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n895_), .A2(new_n286_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n410_), .ZN(G1355gat));
endmodule


