//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n861_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n203_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT79), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(KEYINPUT26), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n213_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n208_), .B(new_n210_), .C1(new_n212_), .C2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT80), .ZN(new_n221_));
  OAI21_X1  g020(.A(G169gat), .B1(new_n221_), .B2(G176gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n219_), .B(new_n222_), .C1(new_n221_), .C2(new_n206_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT81), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n218_), .A2(KEYINPUT81), .A3(new_n223_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n228_), .B(KEYINPUT30), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G71gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231_));
  INV_X1    g030(.A(G113gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G120gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n230_), .A2(new_n236_), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G15gat), .B(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G99gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n242_), .B(new_n244_), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OR3_X1    g045(.A1(new_n238_), .A2(new_n239_), .A3(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n246_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G22gat), .B(G50gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT28), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(G141gat), .A2(G148gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT2), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(KEYINPUT2), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n254_), .A2(new_n257_), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  INV_X1    g060(.A(G155gat), .ZN(new_n262_));
  INV_X1    g061(.A(G162gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n260_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(KEYINPUT1), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n264_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(KEYINPUT83), .A3(new_n264_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n269_), .B(new_n270_), .C1(KEYINPUT1), .C2(new_n261_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n253_), .A2(new_n255_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT84), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT84), .B1(new_n271_), .B2(new_n272_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n265_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n252_), .B1(new_n276_), .B2(KEYINPUT29), .ZN(new_n277_));
  INV_X1    g076(.A(new_n265_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n272_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n281_), .B2(new_n273_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n251_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n277_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT85), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n277_), .A2(KEYINPUT85), .A3(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G197gat), .B(G204gat), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT21), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G211gat), .B(G218gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT86), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n291_), .A2(new_n292_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n301_));
  INV_X1    g100(.A(G228gat), .ZN(new_n302_));
  INV_X1    g101(.A(G233gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n301_), .A2(new_n304_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G78gat), .B(G106gat), .Z(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT87), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n307_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n305_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n310_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n289_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT88), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n308_), .A2(new_n317_), .A3(new_n309_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n309_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT88), .B1(new_n314_), .B2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n285_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n316_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n276_), .A2(new_n236_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n282_), .A2(new_n235_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n325_), .A2(KEYINPUT4), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n325_), .A2(new_n326_), .A3(KEYINPUT4), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT95), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(KEYINPUT95), .A3(KEYINPUT4), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n330_), .B1(new_n336_), .B2(new_n329_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G85gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(G1gat), .B(G29gat), .Z(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n328_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(new_n330_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n205_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n219_), .A2(new_n209_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n211_), .A2(new_n213_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT90), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n203_), .B1(new_n206_), .B2(new_n351_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT91), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n350_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n300_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n298_), .A2(new_n299_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n360_), .A2(new_n369_), .A3(new_n300_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT92), .B1(new_n362_), .B2(new_n359_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(KEYINPUT20), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n366_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT94), .B(G8gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n375_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n366_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n384_), .B1(new_n373_), .B2(new_n366_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n382_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n346_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n345_), .A2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n368_), .A2(new_n374_), .A3(new_n381_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n381_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(KEYINPUT33), .B(new_n343_), .C1(new_n344_), .C2(new_n330_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n327_), .A2(new_n329_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n341_), .B(new_n394_), .C1(new_n336_), .C2(new_n329_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .A4(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n324_), .B1(new_n387_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n381_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n385_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(KEYINPUT27), .C1(new_n400_), .C2(new_n375_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n403_), .A2(new_n323_), .A3(new_n346_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n249_), .B1(new_n397_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n249_), .A2(new_n346_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n324_), .A2(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT96), .B(new_n249_), .C1(new_n397_), .C2(new_n404_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G230gat), .A2(G233gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT10), .B(G99gat), .Z(new_n414_));
  INV_X1    g213(.A(G106gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G85gat), .B(G92gat), .Z(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT9), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n419_));
  INV_X1    g218(.A(G92gat), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT9), .ZN(new_n421_));
  NOR2_X1   g220(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(G85gat), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT6), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n416_), .A2(new_n418_), .A3(new_n423_), .A4(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G71gat), .A2(G78gat), .ZN(new_n430_));
  INV_X1    g229(.A(G71gat), .ZN(new_n431_));
  INV_X1    g230(.A(G78gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G57gat), .B(G64gat), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n430_), .B(new_n433_), .C1(new_n434_), .C2(KEYINPUT11), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT68), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(KEYINPUT11), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n435_), .A2(KEYINPUT68), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(KEYINPUT68), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n439_), .A2(KEYINPUT11), .A3(new_n434_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n428_), .A2(KEYINPUT65), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT66), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT7), .ZN(new_n448_));
  INV_X1    g247(.A(G99gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n415_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n444_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT65), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n425_), .A2(new_n427_), .A3(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n443_), .A2(new_n447_), .A3(new_n452_), .A4(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT67), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n417_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n455_), .B2(new_n417_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT8), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n428_), .A2(new_n450_), .A3(new_n444_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n459_), .A3(new_n417_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n429_), .B(new_n442_), .C1(new_n460_), .C2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT12), .ZN(new_n465_));
  INV_X1    g264(.A(new_n429_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n455_), .A2(new_n417_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT67), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n455_), .A2(new_n456_), .A3(new_n417_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT8), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n466_), .B1(new_n470_), .B2(new_n462_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n471_), .A2(new_n442_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n465_), .A2(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n471_), .A2(KEYINPUT12), .A3(new_n442_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n413_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G120gat), .B(G148gat), .ZN(new_n477_));
  INV_X1    g276(.A(G204gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT5), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(new_n205_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n429_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n442_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(KEYINPUT69), .A3(new_n464_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n413_), .ZN(new_n487_));
  OR3_X1    g286(.A1(new_n471_), .A2(KEYINPUT69), .A3(new_n442_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n476_), .A2(new_n482_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n481_), .B(KEYINPUT70), .Z(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n476_), .B2(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT13), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(KEYINPUT13), .A3(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G1gat), .ZN(new_n499_));
  INV_X1    g298(.A(G8gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT14), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n501_), .A2(KEYINPUT75), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(KEYINPUT75), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G8gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G29gat), .B(G36gat), .ZN(new_n508_));
  INV_X1    g307(.A(G43gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G50gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n511_), .B(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n512_), .B1(new_n514_), .B2(new_n507_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n516_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n507_), .A2(new_n511_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n512_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G169gat), .B(G197gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(G141gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT78), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(new_n232_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n517_), .A2(new_n520_), .A3(new_n525_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n498_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n507_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n484_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G127gat), .B(G155gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT77), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  OR3_X1    g340(.A1(new_n534_), .A2(new_n535_), .A3(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(KEYINPUT17), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT34), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n483_), .B2(new_n514_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n550_));
  OAI221_X1 g349(.A(new_n549_), .B1(KEYINPUT73), .B2(new_n550_), .C1(new_n483_), .C2(new_n511_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n550_), .A2(KEYINPUT73), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n552_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT71), .B(G134gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n263_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT36), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT37), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n561_), .B(KEYINPUT74), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n556_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n566_), .B1(new_n569_), .B2(new_n564_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n545_), .B1(new_n567_), .B2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n412_), .A2(new_n530_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT97), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(new_n499_), .A3(new_n346_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n576_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n412_), .A2(new_n530_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n579_), .A2(new_n565_), .A3(new_n545_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(new_n346_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n577_), .B(new_n578_), .C1(new_n499_), .C2(new_n581_), .ZN(G1324gat));
  AOI21_X1  g381(.A(new_n500_), .B1(new_n580_), .B2(new_n403_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT39), .Z(new_n584_));
  NAND3_X1  g383(.A1(new_n574_), .A2(new_n500_), .A3(new_n403_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT40), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n584_), .A2(KEYINPUT40), .A3(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(G1325gat));
  INV_X1    g389(.A(G15gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n249_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n574_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n580_), .B2(new_n592_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n596_), .A2(KEYINPUT41), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT41), .B1(new_n596_), .B2(new_n597_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n593_), .B1(new_n598_), .B2(new_n599_), .ZN(G1326gat));
  INV_X1    g399(.A(G22gat), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n580_), .B2(new_n324_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT42), .Z(new_n603_));
  NAND3_X1  g402(.A1(new_n574_), .A2(new_n601_), .A3(new_n324_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT99), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n607_), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(G1327gat));
  NAND2_X1  g408(.A1(new_n565_), .A2(new_n545_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT102), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n579_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(G29gat), .B1(new_n613_), .B2(new_n346_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n562_), .A2(new_n564_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(KEYINPUT37), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n570_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n412_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n617_), .A2(KEYINPUT101), .A3(new_n570_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT101), .B1(new_n617_), .B2(new_n570_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n620_), .B1(new_n412_), .B2(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n545_), .B(new_n530_), .C1(new_n619_), .C2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(new_n346_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n626_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(G29gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n614_), .B1(new_n628_), .B2(new_n630_), .ZN(G1328gat));
  INV_X1    g430(.A(G36gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n403_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n627_), .B2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n613_), .A2(new_n632_), .A3(new_n403_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT45), .Z(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n635_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1329gat));
  NAND2_X1  g440(.A1(new_n613_), .A2(new_n592_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n509_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n627_), .A2(new_n592_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n629_), .A2(G43gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT47), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT47), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(new_n643_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1330gat));
  NOR2_X1   g449(.A1(new_n323_), .A2(G50gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT103), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n613_), .A2(new_n652_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n627_), .A2(new_n324_), .A3(new_n629_), .ZN(new_n654_));
  INV_X1    g453(.A(G50gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(G1331gat));
  INV_X1    g455(.A(new_n498_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n529_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n412_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n545_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n617_), .B2(new_n570_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n346_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n660_), .A2(new_n565_), .A3(new_n545_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(new_n346_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n666_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g466(.A(G64gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n665_), .B2(new_n403_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT48), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n663_), .A2(new_n668_), .A3(new_n403_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1333gat));
  AOI21_X1  g471(.A(new_n431_), .B1(new_n665_), .B2(new_n592_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT49), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n663_), .A2(new_n431_), .A3(new_n592_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1334gat));
  AOI21_X1  g475(.A(new_n432_), .B1(new_n665_), .B2(new_n324_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT50), .Z(new_n678_));
  NAND3_X1  g477(.A1(new_n663_), .A2(new_n432_), .A3(new_n324_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1335gat));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n660_), .B2(new_n612_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n412_), .A2(KEYINPUT104), .A3(new_n611_), .A4(new_n659_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n346_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n619_), .A2(new_n624_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n657_), .A2(new_n661_), .A3(new_n658_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT105), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n346_), .A2(G85gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT106), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n689_), .B2(new_n691_), .ZN(G1336gat));
  AOI21_X1  g491(.A(G92gat), .B1(new_n684_), .B2(new_n403_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n419_), .A2(new_n420_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n403_), .B1(new_n422_), .B2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT107), .Z(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n689_), .B2(new_n696_), .ZN(G1337gat));
  NAND2_X1  g496(.A1(new_n689_), .A2(new_n592_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G99gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n684_), .A2(new_n414_), .A3(new_n592_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n700_), .ZN(new_n701_));
  OR2_X1    g500(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n702_));
  NAND2_X1  g501(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n449_), .B1(new_n689_), .B2(new_n592_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n700_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n702_), .B(new_n703_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n701_), .A2(new_n706_), .ZN(G1338gat));
  INV_X1    g506(.A(KEYINPUT52), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n324_), .B(new_n688_), .C1(new_n619_), .C2(new_n624_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G106gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G106gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n709_), .A2(G106gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT110), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(new_n710_), .A3(G106gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(KEYINPUT52), .A3(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n684_), .A2(new_n415_), .A3(new_n324_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT109), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n684_), .A2(new_n720_), .A3(new_n415_), .A4(new_n324_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n713_), .A2(new_n717_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT53), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n713_), .A2(new_n717_), .A3(new_n722_), .A4(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1339gat));
  INV_X1    g526(.A(KEYINPUT54), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n572_), .A2(new_n728_), .A3(new_n529_), .A4(new_n657_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n657_), .A2(new_n529_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT54), .B1(new_n662_), .B2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n475_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n485_), .A2(KEYINPUT12), .A3(new_n464_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n474_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n487_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT111), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n735_), .A2(new_n736_), .A3(new_n739_), .A4(new_n487_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT55), .B(new_n413_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n734_), .A2(new_n738_), .A3(new_n740_), .A4(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n492_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT56), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(KEYINPUT56), .A3(new_n492_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT56), .B1(new_n742_), .B2(new_n492_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n490_), .B1(new_n749_), .B2(KEYINPUT112), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n658_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n515_), .A2(new_n518_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n516_), .B1(new_n519_), .B2(new_n512_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n526_), .A3(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n528_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT113), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n494_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n751_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(KEYINPUT57), .A3(new_n616_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n616_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n745_), .A2(new_n765_), .A3(new_n747_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n742_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n492_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(new_n756_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n768_), .A3(new_n491_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n766_), .A2(new_n768_), .A3(KEYINPUT58), .A4(new_n491_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n618_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n565_), .B1(new_n751_), .B2(new_n757_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n761_), .A2(new_n764_), .A3(new_n773_), .A4(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n732_), .B1(new_n776_), .B2(new_n545_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n592_), .A2(new_n346_), .A3(new_n409_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT116), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  INV_X1    g579(.A(new_n778_), .ZN(new_n781_));
  AND4_X1   g580(.A1(KEYINPUT115), .A2(new_n758_), .A3(KEYINPUT57), .A4(new_n616_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT115), .B1(new_n774_), .B2(KEYINPUT57), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n771_), .A2(new_n772_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n785_), .A2(new_n618_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n661_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n780_), .B(new_n781_), .C1(new_n787_), .C2(new_n732_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n779_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(G113gat), .B1(new_n789_), .B2(new_n658_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n787_), .B2(new_n732_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n792_), .B(new_n793_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n777_), .B2(KEYINPUT117), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n777_), .A2(new_n778_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n529_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n790_), .B1(new_n798_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g598(.A(new_n234_), .B1(new_n657_), .B2(KEYINPUT60), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n789_), .B(new_n800_), .C1(KEYINPUT60), .C2(new_n234_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n657_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n234_), .ZN(G1341gat));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  INV_X1    g603(.A(G127gat), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n545_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G127gat), .B1(new_n789_), .B2(new_n661_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n804_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n776_), .A2(new_n545_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n732_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n780_), .B1(new_n813_), .B2(new_n781_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n777_), .A2(KEYINPUT116), .A3(new_n778_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n661_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n805_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n795_), .A2(new_n796_), .ZN(new_n818_));
  AOI221_X4 g617(.A(new_n778_), .B1(KEYINPUT117), .B2(new_n793_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n806_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(KEYINPUT118), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n810_), .A2(new_n821_), .ZN(G1342gat));
  AOI21_X1  g621(.A(G134gat), .B1(new_n789_), .B2(new_n565_), .ZN(new_n823_));
  INV_X1    g622(.A(G134gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n825_), .B2(new_n618_), .ZN(G1343gat));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  INV_X1    g626(.A(new_n346_), .ZN(new_n828_));
  NOR4_X1   g627(.A1(new_n592_), .A2(new_n828_), .A3(new_n323_), .A4(new_n403_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n813_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n829_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT119), .B1(new_n777_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n658_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n498_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g636(.A1(new_n833_), .A2(new_n661_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(new_n262_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT120), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n838_), .B(new_n841_), .ZN(G1346gat));
  AND3_X1   g641(.A1(new_n833_), .A2(G162gat), .A3(new_n623_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n616_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n263_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT122), .B1(new_n844_), .B2(G162gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n843_), .B1(new_n847_), .B2(new_n848_), .ZN(G1347gat));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n777_), .A2(new_n346_), .A3(new_n249_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n633_), .A2(new_n324_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n529_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n850_), .B1(new_n854_), .B2(new_n204_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n347_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT62), .B(G169gat), .C1(new_n853_), .C2(new_n529_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(G1348gat));
  NOR2_X1   g657(.A1(new_n853_), .A2(new_n657_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(new_n205_), .ZN(G1349gat));
  NAND3_X1  g659(.A1(new_n851_), .A2(new_n661_), .A3(new_n852_), .ZN(new_n861_));
  MUX2_X1   g660(.A(new_n213_), .B(G183gat), .S(new_n861_), .Z(G1350gat));
  AND4_X1   g661(.A1(new_n408_), .A2(new_n813_), .A3(new_n618_), .A4(new_n852_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n565_), .A2(new_n211_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT123), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n215_), .A2(new_n863_), .B1(new_n853_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT124), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868_));
  OAI221_X1 g667(.A(new_n868_), .B1(new_n853_), .B2(new_n865_), .C1(new_n215_), .C2(new_n863_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1351gat));
  NOR3_X1   g669(.A1(new_n592_), .A2(new_n323_), .A3(new_n633_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n813_), .A2(new_n828_), .A3(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n529_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT125), .B(G197gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1352gat));
  NOR2_X1   g674(.A1(new_n872_), .A2(new_n657_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n478_), .ZN(G1353gat));
  NOR2_X1   g676(.A1(new_n777_), .A2(new_n346_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n878_), .A2(new_n661_), .A3(new_n871_), .A4(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n881_), .A2(KEYINPUT126), .A3(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT126), .B1(new_n881_), .B2(new_n883_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n879_), .B1(new_n872_), .B2(new_n545_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT127), .B(new_n879_), .C1(new_n872_), .C2(new_n545_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n884_), .A2(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1354gat));
  INV_X1    g689(.A(G218gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n872_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n878_), .A2(new_n565_), .A3(new_n871_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n892_), .A2(new_n618_), .B1(new_n893_), .B2(new_n891_), .ZN(G1355gat));
endmodule


