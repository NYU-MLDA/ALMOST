//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G225gat), .A2(G233gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207_));
  INV_X1    g006(.A(G134gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G127gat), .ZN(new_n209_));
  INV_X1    g008(.A(G127gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G134gat), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT78), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT78), .B1(new_n209_), .B2(new_n211_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G113gat), .B(G120gat), .Z(new_n214_));
  NOR3_X1   g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G113gat), .B(G120gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT78), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n210_), .A2(G134gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n208_), .A2(G127gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT78), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n207_), .B1(new_n215_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n214_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n221_), .A3(new_n216_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT79), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n228_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(KEYINPUT1), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT81), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(new_n229_), .B2(KEYINPUT1), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n232_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G141gat), .ZN(new_n238_));
  INV_X1    g037(.A(G148gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G141gat), .A2(G148gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT82), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT3), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n248_), .A2(new_n238_), .A3(new_n239_), .A4(KEYINPUT82), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT83), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n230_), .A2(new_n228_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n242_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n227_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT4), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n224_), .A2(new_n225_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT98), .B1(new_n255_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n240_), .A2(new_n241_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n233_), .B(KEYINPUT81), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(new_n232_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n250_), .A2(new_n252_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT83), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT98), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n225_), .A4(new_n224_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n227_), .A2(new_n255_), .A3(KEYINPUT97), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT97), .B1(new_n227_), .B2(new_n255_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n260_), .B(new_n269_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  AOI211_X1 g071(.A(new_n206_), .B(new_n258_), .C1(new_n272_), .C2(KEYINPUT4), .ZN(new_n273_));
  INV_X1    g072(.A(new_n206_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n269_), .A2(new_n260_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT97), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n256_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n227_), .A2(new_n255_), .A3(KEYINPUT97), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n274_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n205_), .B1(new_n273_), .B2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n258_), .B1(new_n272_), .B2(KEYINPUT4), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n274_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n205_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n280_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G8gat), .B(G36gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT18), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G64gat), .B(G92gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT19), .Z(new_n294_));
  INV_X1    g093(.A(G197gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(G204gat), .ZN(new_n296_));
  INV_X1    g095(.A(G204gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(G197gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT21), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G211gat), .B(G218gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT86), .B1(new_n295_), .B2(G204gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT86), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(new_n297_), .A3(G197gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n301_), .B(new_n303_), .C1(G197gat), .C2(new_n297_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n299_), .B(new_n300_), .C1(new_n304_), .C2(KEYINPUT21), .ZN(new_n305_));
  INV_X1    g104(.A(new_n300_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(KEYINPUT21), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT95), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(KEYINPUT95), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT96), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT96), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n313_), .A2(new_n319_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT23), .ZN(new_n322_));
  OR2_X1    g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G169gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n312_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n330_), .A2(KEYINPUT24), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(KEYINPUT24), .A3(new_n314_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n328_), .A2(new_n322_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n310_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT22), .B1(new_n337_), .B2(new_n329_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n329_), .A2(KEYINPUT22), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n312_), .B(new_n338_), .C1(new_n339_), .C2(new_n337_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n324_), .A2(new_n314_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n332_), .B(KEYINPUT76), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n328_), .A2(new_n322_), .A3(new_n331_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n336_), .B1(new_n344_), .B2(new_n308_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n294_), .B1(new_n335_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT20), .B1(new_n344_), .B2(new_n308_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n333_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n333_), .A2(new_n348_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n325_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n347_), .B1(new_n308_), .B2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n294_), .B(KEYINPUT93), .Z(new_n353_));
  AND2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n292_), .B1(new_n346_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n292_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n308_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n357_), .A2(new_n325_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n345_), .A3(new_n294_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n356_), .B(new_n359_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n360_), .A2(KEYINPUT27), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n351_), .A2(new_n308_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n347_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n353_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n359_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n292_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n367_), .A2(new_n360_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n362_), .B1(KEYINPUT27), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT88), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n267_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n255_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n310_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n267_), .B2(new_n372_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(KEYINPUT87), .B(new_n378_), .C1(new_n267_), .C2(new_n372_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n375_), .A2(new_n377_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G78gat), .B(G106gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT90), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT91), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G22gat), .B(G50gat), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n242_), .B(new_n372_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT84), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n265_), .A2(new_n266_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT84), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n372_), .A4(new_n242_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n390_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n388_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n267_), .B2(new_n372_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n389_), .A2(KEYINPUT84), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n394_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n390_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n387_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT92), .B1(new_n386_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n375_), .A2(new_n377_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n381_), .A2(new_n382_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n385_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n398_), .A2(new_n403_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT92), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n406_), .A2(new_n407_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(new_n385_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n405_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n405_), .B2(new_n413_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n288_), .B(new_n370_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(new_n359_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n346_), .A2(new_n354_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n419_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n272_), .A2(KEYINPUT4), .ZN(new_n424_));
  INV_X1    g223(.A(new_n258_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n274_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n284_), .B1(new_n272_), .B2(new_n206_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n368_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n280_), .B1(new_n282_), .B2(new_n274_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT99), .B1(new_n429_), .B2(new_n284_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n430_), .B2(KEYINPUT33), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n281_), .A2(KEYINPUT99), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n423_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n383_), .B(new_n385_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n386_), .A2(KEYINPUT92), .A3(new_n404_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n412_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n405_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n418_), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(G15gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT30), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n344_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(new_n227_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G43gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT31), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n447_), .B(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n452_), .B(KEYINPUT80), .Z(new_n453_));
  NOR2_X1   g252(.A1(new_n416_), .A2(new_n417_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n281_), .A2(new_n286_), .A3(new_n452_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(KEYINPUT100), .A3(new_n370_), .A4(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n438_), .A2(new_n455_), .A3(new_n370_), .A4(new_n439_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT100), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n441_), .A2(new_n453_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n461_));
  INV_X1    g260(.A(G1gat), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G8gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n465_), .B(new_n466_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n470_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n473_), .A2(new_n474_), .A3(KEYINPUT73), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n476_), .A2(G229gat), .A3(G233gat), .A4(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n470_), .B(KEYINPUT15), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT74), .Z(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n471_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G169gat), .B(G197gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n478_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT75), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT75), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n484_), .A2(new_n492_), .A3(new_n488_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n460_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G120gat), .B(G148gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT5), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G176gat), .B(G204gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT65), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G230gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n504_), .A2(KEYINPUT64), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(KEYINPUT64), .ZN(new_n506_));
  OR3_X1    g305(.A1(new_n505_), .A2(new_n506_), .A3(KEYINPUT11), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT11), .B1(new_n505_), .B2(new_n506_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n508_), .A2(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G85gat), .B(G92gat), .Z(new_n514_));
  NOR2_X1   g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n514_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT8), .ZN(new_n522_));
  INV_X1    g321(.A(new_n520_), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT10), .B(G99gat), .Z(new_n524_));
  INV_X1    g323(.A(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n514_), .A2(KEYINPUT9), .ZN(new_n527_));
  INV_X1    g326(.A(G85gat), .ZN(new_n528_));
  INV_X1    g327(.A(G92gat), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT9), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n523_), .A2(new_n526_), .A3(new_n527_), .A4(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n522_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n513_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n512_), .A2(new_n531_), .A3(new_n522_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(KEYINPUT12), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n513_), .A2(new_n536_), .A3(new_n532_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n503_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n502_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n501_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n538_), .A2(new_n539_), .A3(new_n501_), .ZN(new_n543_));
  OR3_X1    g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n532_), .A2(new_n479_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n522_), .A2(new_n470_), .A3(new_n531_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT67), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT66), .B(KEYINPUT34), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n549_), .A2(new_n550_), .A3(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n554_), .A2(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n563_));
  INV_X1    g362(.A(new_n558_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n549_), .A2(new_n564_), .A3(new_n550_), .A4(new_n556_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n559_), .A2(new_n565_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n562_), .B(KEYINPUT36), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n548_), .B(new_n566_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n566_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n571_), .A2(new_n572_), .A3(KEYINPUT69), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n570_), .B1(new_n573_), .B2(new_n548_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT37), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT70), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT69), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n577_), .B(new_n566_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT37), .B1(new_n578_), .B2(KEYINPUT68), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(new_n576_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT37), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(KEYINPUT68), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(new_n570_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT70), .B1(new_n584_), .B2(new_n579_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n512_), .A2(new_n467_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(G231gat), .ZN(new_n590_));
  INV_X1    g389(.A(G233gat), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n473_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n588_), .B2(new_n594_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT17), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n596_), .A2(new_n597_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n603_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n596_), .A2(new_n597_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT72), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT72), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n596_), .A2(new_n597_), .A3(new_n604_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n596_), .A2(new_n597_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n604_), .A2(new_n606_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n609_), .B(new_n610_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n587_), .A2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n495_), .A2(new_n547_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n462_), .A3(new_n287_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n571_), .A2(new_n572_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n460_), .A2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n546_), .A2(new_n494_), .A3(new_n614_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n288_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n617_), .A2(new_n618_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n619_), .A2(new_n624_), .A3(new_n625_), .ZN(G1324gat));
  NAND3_X1  g425(.A1(new_n616_), .A2(new_n463_), .A3(new_n369_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n623_), .A2(new_n370_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n463_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT101), .B1(new_n623_), .B2(new_n370_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n627_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(G1325gat));
  OAI21_X1  g436(.A(G15gat), .B1(new_n623_), .B2(new_n453_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT41), .Z(new_n639_));
  INV_X1    g438(.A(new_n453_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n616_), .A2(new_n443_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(G1326gat));
  OAI21_X1  g441(.A(G22gat), .B1(new_n623_), .B2(new_n454_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(G22gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n616_), .A2(new_n646_), .A3(new_n440_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1327gat));
  OAI21_X1  g447(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n586_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n430_), .A2(KEYINPUT33), .ZN(new_n651_));
  INV_X1    g450(.A(new_n428_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n433_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n423_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n454_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n640_), .B1(new_n656_), .B2(new_n418_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n457_), .B(KEYINPUT100), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n650_), .B(new_n587_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n649_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n494_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n547_), .A2(new_n661_), .A3(new_n614_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(KEYINPUT44), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT104), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n662_), .B1(new_n649_), .B2(new_n659_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n441_), .A2(new_n453_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n456_), .A2(new_n459_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n650_), .B1(new_n672_), .B2(new_n587_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n460_), .A2(KEYINPUT43), .A3(new_n586_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n663_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(KEYINPUT103), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(new_n666_), .B2(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n669_), .A2(new_n680_), .A3(new_n287_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G29gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n614_), .A2(new_n620_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT105), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(new_n546_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n495_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n288_), .A2(G29gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT106), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n682_), .B1(new_n686_), .B2(new_n688_), .ZN(G1328gat));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n669_), .A2(new_n680_), .A3(new_n369_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n370_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n686_), .B2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n495_), .A2(new_n685_), .A3(new_n696_), .A4(new_n698_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n690_), .A2(new_n691_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n693_), .B1(new_n695_), .B2(new_n705_), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n692_), .B(new_n704_), .C1(new_n694_), .C2(G36gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1329gat));
  NAND4_X1  g507(.A1(new_n669_), .A2(new_n680_), .A3(G43gat), .A4(new_n452_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n449_), .B1(new_n686_), .B2(new_n453_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT47), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n713_), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1330gat));
  NAND3_X1  g514(.A1(new_n669_), .A2(new_n680_), .A3(new_n440_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(G50gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G50gat), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n454_), .A2(G50gat), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT110), .ZN(new_n721_));
  OAI22_X1  g520(.A1(new_n718_), .A2(new_n719_), .B1(new_n686_), .B2(new_n721_), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n615_), .A2(new_n546_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT111), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n672_), .A3(new_n494_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT112), .ZN(new_n726_));
  INV_X1    g525(.A(G57gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n287_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n547_), .A2(new_n661_), .A3(new_n614_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n621_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n288_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(G1332gat));
  INV_X1    g532(.A(G64gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n726_), .A2(new_n734_), .A3(new_n369_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n730_), .B2(new_n369_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT48), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n726_), .A2(new_n739_), .A3(new_n640_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n730_), .B2(new_n640_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT49), .Z(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1334gat));
  INV_X1    g542(.A(G78gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n726_), .A2(new_n744_), .A3(new_n440_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n730_), .B2(new_n440_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT50), .Z(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1335gat));
  INV_X1    g547(.A(new_n614_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n547_), .A2(new_n661_), .A3(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n660_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n288_), .ZN(new_n753_));
  NOR4_X1   g552(.A1(new_n460_), .A2(new_n661_), .A3(new_n547_), .A4(new_n684_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n528_), .A3(new_n287_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT113), .Z(G1336gat));
  AOI21_X1  g556(.A(G92gat), .B1(new_n754_), .B2(new_n369_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n369_), .A2(G92gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT114), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n751_), .B2(new_n760_), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n752_), .B2(new_n453_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n452_), .A2(new_n524_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n754_), .A2(new_n763_), .B1(new_n764_), .B2(KEYINPUT51), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(KEYINPUT51), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n766_), .B(new_n767_), .Z(G1338gat));
  NAND3_X1  g567(.A1(new_n754_), .A2(new_n525_), .A3(new_n440_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n751_), .A2(new_n440_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G106gat), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT52), .B(new_n525_), .C1(new_n751_), .C2(new_n440_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XOR2_X1   g573(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n775_));
  XNOR2_X1  g574(.A(new_n774_), .B(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT124), .ZN(new_n777_));
  INV_X1    g576(.A(G113gat), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT123), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n454_), .A2(new_n287_), .A3(new_n370_), .A4(new_n452_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT121), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(KEYINPUT59), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n535_), .A2(new_n537_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n502_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n535_), .A2(new_n503_), .A3(new_n537_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(KEYINPUT55), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n500_), .B1(new_n538_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n538_), .A2(new_n539_), .A3(new_n499_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n482_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n487_), .B1(new_n480_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n476_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n490_), .A2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n792_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n791_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n788_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT58), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n800_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n791_), .A4(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n792_), .A2(new_n494_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n787_), .A2(new_n790_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n541_), .A2(new_n543_), .ZN(new_n812_));
  OAI22_X1  g611(.A1(new_n810_), .A2(new_n811_), .B1(new_n812_), .B2(new_n797_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n620_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n814_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n806_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT122), .B1(new_n819_), .B2(new_n614_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT117), .B1(new_n614_), .B2(new_n661_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n608_), .A2(new_n613_), .A3(new_n822_), .A4(new_n494_), .ZN(new_n823_));
  AND4_X1   g622(.A1(new_n544_), .A2(new_n821_), .A3(new_n545_), .A4(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n576_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n584_), .A2(KEYINPUT70), .A3(new_n579_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(KEYINPUT54), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(KEYINPUT54), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n586_), .A2(new_n828_), .A3(KEYINPUT54), .A4(new_n824_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n820_), .A2(new_n834_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n819_), .A2(KEYINPUT122), .A3(new_n614_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n779_), .B(new_n783_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n836_), .A2(new_n820_), .A3(new_n834_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n783_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT123), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  INV_X1    g640(.A(new_n818_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n814_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n806_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n805_), .A2(new_n581_), .A3(new_n585_), .A4(KEYINPUT120), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n614_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n832_), .A2(new_n833_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n841_), .B1(new_n851_), .B2(new_n781_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n837_), .B1(new_n840_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n778_), .B1(new_n853_), .B2(new_n661_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n834_), .B1(new_n614_), .B2(new_n848_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n782_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n778_), .A3(new_n661_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n777_), .B1(new_n854_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n783_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT59), .B1(new_n855_), .B2(new_n782_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(KEYINPUT123), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n494_), .B1(new_n862_), .B2(new_n837_), .ZN(new_n863_));
  OAI211_X1 g662(.A(KEYINPUT124), .B(new_n857_), .C1(new_n863_), .C2(new_n778_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(G1340gat));
  INV_X1    g664(.A(G120gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n547_), .B2(KEYINPUT60), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n856_), .B(new_n867_), .C1(KEYINPUT60), .C2(new_n866_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n547_), .B1(new_n862_), .B2(new_n837_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n866_), .ZN(G1341gat));
  NAND3_X1  g669(.A1(new_n856_), .A2(new_n210_), .A3(new_n749_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n614_), .B1(new_n862_), .B2(new_n837_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n210_), .ZN(G1342gat));
  NAND3_X1  g672(.A1(new_n856_), .A2(new_n208_), .A3(new_n620_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n586_), .B1(new_n862_), .B2(new_n837_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n208_), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n640_), .A2(new_n288_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n851_), .A2(new_n440_), .A3(new_n370_), .A4(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n494_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n238_), .ZN(G1344gat));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n547_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n239_), .ZN(G1345gat));
  NOR2_X1   g681(.A1(new_n878_), .A2(new_n614_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT61), .B(G155gat), .Z(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  OAI21_X1  g684(.A(G162gat), .B1(new_n878_), .B2(new_n586_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n814_), .A2(G162gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n878_), .B2(new_n887_), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n838_), .A2(new_n440_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n453_), .A2(new_n287_), .A3(new_n370_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891_), .B2(new_n494_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n893_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n891_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n311_), .A3(new_n661_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n895_), .A3(new_n897_), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n896_), .B2(new_n546_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n855_), .A2(new_n440_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n890_), .A2(G176gat), .A3(new_n546_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  NAND2_X1  g701(.A1(new_n890_), .A2(new_n749_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G183gat), .B1(new_n900_), .B2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n326_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n889_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n891_), .B2(new_n586_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n620_), .A2(new_n327_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT126), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n891_), .B2(new_n912_), .ZN(G1351gat));
  NOR4_X1   g712(.A1(new_n640_), .A2(new_n454_), .A3(new_n287_), .A4(new_n370_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n851_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n494_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n295_), .ZN(G1352gat));
  INV_X1    g716(.A(new_n915_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n918_), .B(new_n546_), .C1(KEYINPUT127), .C2(new_n297_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n297_), .A2(KEYINPUT127), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1353gat));
  NOR2_X1   g720(.A1(new_n915_), .A2(new_n614_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AND2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n922_), .B2(new_n923_), .ZN(G1354gat));
  OR3_X1    g725(.A1(new_n915_), .A2(G218gat), .A3(new_n814_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G218gat), .B1(new_n915_), .B2(new_n586_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1355gat));
endmodule


