//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G155gat), .ZN(new_n206_));
  INV_X1    g005(.A(G162gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  AOI211_X1 g020(.A(new_n208_), .B(new_n209_), .C1(new_n218_), .C2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G141gat), .B(G148gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n208_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT1), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n209_), .B1(new_n208_), .B2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n223_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n205_), .B1(new_n222_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n221_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n209_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n224_), .A3(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n225_), .A2(new_n227_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n232_), .B(new_n204_), .C1(new_n233_), .C2(new_n223_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n229_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n229_), .A2(new_n234_), .A3(KEYINPUT4), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n235_), .B(KEYINPUT91), .Z(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n229_), .B2(KEYINPUT4), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n236_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G1gat), .B(G29gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G85gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT0), .B(G57gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n236_), .B(new_n246_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n204_), .B(KEYINPUT31), .Z(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G99gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(G43gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT78), .B(G15gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G227gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT22), .B(G169gat), .ZN(new_n259_));
  INV_X1    g058(.A(G176gat), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT23), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT76), .B(G183gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(G190gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n261_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT24), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n258_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n269_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n263_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n272_), .B2(KEYINPUT77), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n263_), .A2(new_n271_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n276_), .B1(new_n265_), .B2(KEYINPUT25), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT26), .B(G190gat), .Z(new_n278_));
  OAI22_X1  g077(.A1(new_n274_), .A2(new_n275_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n267_), .B1(new_n273_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT30), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT79), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n256_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n256_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n250_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n287_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n250_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n285_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n249_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT97), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT27), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  NAND3_X1  g094(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G211gat), .B(G218gat), .Z(new_n300_));
  OR2_X1    g099(.A1(G197gat), .A2(G204gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT82), .B(G204gat), .ZN(new_n302_));
  INV_X1    g101(.A(G197gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT21), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n302_), .A2(G197gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n303_), .A2(G204gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT21), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(KEYINPUT84), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n300_), .A2(KEYINPUT83), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n313_), .B(new_n301_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n305_), .B1(new_n300_), .B2(KEYINPUT83), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  AOI211_X1 g116(.A(new_n295_), .B(new_n299_), .C1(new_n280_), .C2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT25), .B(G183gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT88), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n270_), .B(new_n272_), .C1(new_n320_), .C2(new_n278_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n261_), .B1(new_n264_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT89), .B1(new_n324_), .B2(new_n317_), .ZN(new_n325_));
  OR3_X1    g124(.A1(new_n324_), .A2(new_n317_), .A3(KEYINPUT89), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n318_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n299_), .B(KEYINPUT87), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n280_), .A2(new_n317_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n295_), .B1(new_n324_), .B2(new_n317_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT18), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G64gat), .B(G92gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n327_), .A2(new_n332_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n332_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n318_), .A2(new_n326_), .A3(new_n325_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n294_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n324_), .A2(new_n317_), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n280_), .B2(new_n317_), .ZN(new_n345_));
  AOI211_X1 g144(.A(new_n298_), .B(new_n297_), .C1(new_n343_), .C2(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n330_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n336_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n339_), .A2(new_n340_), .A3(new_n338_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT27), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n342_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT85), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT29), .B1(new_n222_), .B2(new_n228_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n317_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(KEYINPUT81), .A2(G233gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(G228gat), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n317_), .A3(new_n359_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n353_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n353_), .A3(new_n362_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n222_), .A2(KEYINPUT29), .A3(new_n228_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G22gat), .B(G50gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT28), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n367_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT86), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n370_), .B1(new_n363_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n366_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n364_), .A2(new_n371_), .A3(new_n365_), .A4(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n293_), .B1(new_n351_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n377_), .A2(new_n342_), .A3(KEYINPUT97), .A4(new_n350_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n292_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n351_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n377_), .A2(new_n248_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n336_), .A2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n384_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n248_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n384_), .B(KEYINPUT94), .Z(new_n387_));
  INV_X1    g186(.A(KEYINPUT95), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT95), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n386_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n337_), .A2(new_n341_), .A3(KEYINPUT90), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n336_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(new_n349_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n229_), .A2(new_n234_), .A3(new_n238_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n244_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n399_), .A2(KEYINPUT93), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(KEYINPUT93), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n235_), .B1(new_n229_), .B2(KEYINPUT4), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n400_), .B(new_n401_), .C1(new_n237_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n247_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT33), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT92), .B1(new_n404_), .B2(KEYINPUT33), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT92), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n247_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n392_), .B1(new_n397_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n382_), .B1(new_n412_), .B2(new_n375_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n288_), .A2(new_n291_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n379_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G29gat), .B(G36gat), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n416_), .A2(KEYINPUT70), .ZN(new_n417_));
  INV_X1    g216(.A(G36gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G29gat), .ZN(new_n419_));
  INV_X1    g218(.A(G29gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G36gat), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n419_), .A2(new_n421_), .A3(KEYINPUT70), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G43gat), .B(G50gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n416_), .A2(KEYINPUT70), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n422_), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n429_));
  AND3_X1   g228(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G1gat), .ZN(new_n433_));
  INV_X1    g232(.A(G8gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT74), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT74), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n437_), .B(KEYINPUT14), .C1(new_n433_), .C2(new_n434_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G1gat), .B(G8gat), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n441_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n432_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n444_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n425_), .A2(new_n428_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n446_), .A2(new_n447_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n447_), .A2(new_n443_), .A3(new_n442_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n450_), .B1(new_n453_), .B2(new_n449_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G113gat), .B(G141gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G169gat), .B(G197gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n450_), .B(new_n457_), .C1(new_n453_), .C2(new_n449_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n415_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G190gat), .B(G218gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G134gat), .B(G162gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT36), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467_));
  INV_X1    g266(.A(G99gat), .ZN(new_n468_));
  INV_X1    g267(.A(G106gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(KEYINPUT65), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n474_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(KEYINPUT65), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n473_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n472_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G85gat), .B(G92gat), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT8), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n470_), .A2(new_n471_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n480_), .A2(new_n481_), .A3(new_n473_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n473_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n484_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT68), .ZN(new_n494_));
  INV_X1    g293(.A(G85gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT64), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT64), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G85gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G92gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n501_));
  INV_X1    g300(.A(G92gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n495_), .A2(new_n502_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n500_), .A2(new_n501_), .B1(KEYINPUT9), .B2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n469_), .A3(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n494_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n505_), .A2(new_n506_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n479_), .A2(new_n482_), .B1(new_n510_), .B2(new_n469_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n503_), .A2(KEYINPUT9), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n502_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n501_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(KEYINPUT68), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n493_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n432_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n486_), .A2(new_n492_), .B1(new_n515_), .B2(new_n511_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n447_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT34), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n518_), .A2(new_n520_), .A3(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n524_), .A2(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n518_), .A2(new_n530_), .A3(new_n520_), .A4(new_n526_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n466_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n465_), .A2(KEYINPUT36), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n533_), .A3(new_n531_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT73), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n529_), .A2(KEYINPUT73), .A3(new_n533_), .A4(new_n531_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n532_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(KEYINPUT37), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540_));
  AOI211_X1 g339(.A(new_n540_), .B(new_n532_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  XOR2_X1   g343(.A(G71gat), .B(G78gat), .Z(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n444_), .B(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G127gat), .B(G155gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT16), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT17), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT75), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT75), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561_));
  OR3_X1    g360(.A1(new_n552_), .A2(new_n561_), .A3(new_n556_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n542_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT5), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n511_), .A2(new_n515_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n483_), .A2(KEYINPUT8), .A3(new_n485_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n491_), .B1(new_n490_), .B2(new_n484_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n571_), .B(new_n549_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n493_), .A2(KEYINPUT66), .A3(new_n571_), .A4(new_n549_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(KEYINPUT67), .A3(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n549_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT67), .B1(new_n576_), .B2(new_n577_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n570_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(new_n519_), .B2(new_n549_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n570_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n519_), .B2(new_n549_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n546_), .B(KEYINPUT12), .C1(new_n547_), .C2(new_n548_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n572_), .A2(new_n573_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n509_), .A2(new_n516_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n587_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT69), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n587_), .A2(new_n589_), .A3(new_n594_), .A4(KEYINPUT69), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n569_), .B1(new_n585_), .B2(new_n599_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n581_), .A2(new_n586_), .B1(new_n517_), .B2(new_n591_), .ZN(new_n601_));
  AOI21_X1  g400(.A(KEYINPUT69), .B1(new_n601_), .B2(new_n589_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n598_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n578_), .A2(new_n581_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n588_), .B1(new_n605_), .B2(new_n583_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n569_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n600_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT13), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n600_), .A2(KEYINPUT13), .A3(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n565_), .A2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n462_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT98), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n433_), .A3(new_n248_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n415_), .A2(new_n563_), .A3(new_n538_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n613_), .A2(new_n461_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n249_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n617_), .A2(new_n618_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n619_), .A2(new_n624_), .A3(new_n625_), .ZN(G1324gat));
  NOR2_X1   g425(.A1(new_n380_), .A2(G8gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n616_), .A2(new_n627_), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT39), .B(new_n434_), .C1(new_n622_), .C2(new_n351_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n622_), .A2(new_n351_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n631_), .B2(G8gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n628_), .B(KEYINPUT40), .C1(new_n629_), .C2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1325gat));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n462_), .A2(new_n614_), .ZN(new_n639_));
  OR4_X1    g438(.A1(new_n638_), .A2(new_n639_), .A3(G15gat), .A4(new_n414_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n414_), .A2(G15gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n644_));
  INV_X1    g443(.A(new_n414_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n622_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n646_), .B2(G15gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n644_), .A3(G15gat), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n643_), .A2(KEYINPUT100), .A3(new_n648_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n652_), .B2(new_n647_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(G22gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n615_), .A2(new_n655_), .A3(new_n375_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n622_), .A2(new_n375_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G22gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT42), .B(new_n655_), .C1(new_n622_), .C2(new_n375_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT101), .B(new_n656_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1327gat));
  NAND2_X1  g464(.A1(new_n563_), .A2(new_n538_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n613_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n462_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n248_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n613_), .A2(new_n564_), .A3(new_n461_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  INV_X1    g471(.A(new_n392_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n406_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT90), .B1(new_n337_), .B2(new_n341_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n407_), .A2(new_n410_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n395_), .A2(new_n394_), .A3(new_n349_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n375_), .B1(new_n673_), .B2(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n351_), .A2(new_n377_), .A3(new_n248_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n414_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n379_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n542_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n672_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT43), .B(new_n542_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n671_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n687_), .A2(G29gat), .A3(new_n248_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n415_), .B2(new_n542_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n683_), .A2(new_n672_), .A3(new_n684_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n691_), .B2(new_n671_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n670_), .B1(new_n688_), .B2(new_n693_), .ZN(G1328gat));
  XNOR2_X1  g493(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n687_), .A2(new_n351_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G36gat), .B1(new_n696_), .B2(new_n692_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n462_), .A2(new_n418_), .A3(new_n351_), .A4(new_n667_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n695_), .B1(new_n701_), .B2(KEYINPUT103), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703_));
  INV_X1    g502(.A(new_n695_), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n703_), .B(new_n704_), .C1(new_n697_), .C2(new_n700_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n702_), .A2(new_n705_), .ZN(G1329gat));
  NAND3_X1  g505(.A1(new_n687_), .A2(G43gat), .A3(new_n645_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n668_), .A2(new_n414_), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n707_), .A2(new_n692_), .B1(G43gat), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n687_), .A2(G50gat), .A3(new_n375_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n668_), .A2(new_n377_), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n711_), .A2(new_n692_), .B1(G50gat), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT105), .Z(G1331gat));
  INV_X1    g513(.A(new_n461_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n613_), .ZN(new_n716_));
  NOR4_X1   g515(.A1(new_n415_), .A2(new_n715_), .A3(new_n716_), .A4(new_n565_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n248_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n620_), .A2(new_n461_), .A3(new_n613_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(new_n248_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n721_), .B2(new_n718_), .ZN(G1332gat));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n720_), .B2(new_n351_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT48), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n717_), .A2(new_n723_), .A3(new_n351_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n717_), .A2(new_n728_), .A3(new_n645_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT49), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n720_), .A2(new_n645_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G71gat), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT49), .B(new_n728_), .C1(new_n720_), .C2(new_n645_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT106), .B(new_n729_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n720_), .B2(new_n375_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT50), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n717_), .A2(new_n739_), .A3(new_n375_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1335gat));
  NOR3_X1   g542(.A1(new_n716_), .A2(new_n715_), .A3(new_n564_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n691_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n248_), .A3(new_n499_), .ZN(new_n746_));
  NOR4_X1   g545(.A1(new_n415_), .A2(new_n715_), .A3(new_n716_), .A4(new_n666_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n248_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(G85gat), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT107), .ZN(G1336gat));
  AOI21_X1  g549(.A(G92gat), .B1(new_n747_), .B2(new_n351_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT108), .Z(new_n752_));
  NOR2_X1   g551(.A1(new_n380_), .A2(new_n502_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n745_), .B2(new_n753_), .ZN(G1337gat));
  NAND3_X1  g553(.A1(new_n747_), .A2(new_n645_), .A3(new_n510_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n691_), .A2(new_n645_), .A3(new_n744_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n756_), .A2(KEYINPUT109), .A3(G99gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT109), .B1(new_n756_), .B2(G99gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n747_), .A2(new_n469_), .A3(new_n375_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n691_), .A2(new_n375_), .A3(new_n744_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G106gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G106gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g566(.A(new_n414_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n445_), .A2(G229gat), .A3(G233gat), .A4(new_n448_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n449_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n458_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT113), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n769_), .A2(new_n770_), .A3(new_n773_), .A4(new_n458_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n460_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n607_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT114), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n609_), .A2(new_n781_), .A3(new_n776_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n576_), .A2(new_n577_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT111), .B1(new_n783_), .B2(new_n601_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n587_), .A2(new_n594_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n576_), .A2(new_n577_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n588_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n597_), .A2(new_n790_), .A3(new_n598_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n595_), .A2(new_n790_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(KEYINPUT112), .A2(KEYINPUT56), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n569_), .A3(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n777_), .A2(new_n461_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n794_), .B2(new_n569_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n780_), .B(new_n782_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n538_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n597_), .A2(new_n790_), .A3(new_n598_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n783_), .A2(new_n601_), .A3(KEYINPUT111), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n787_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n570_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n804_), .A2(new_n807_), .A3(new_n792_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n607_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n794_), .A2(new_n810_), .A3(new_n569_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n777_), .A2(new_n775_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n542_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n809_), .A2(KEYINPUT58), .A3(new_n811_), .A4(new_n812_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n802_), .A2(new_n803_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n781_), .B1(new_n609_), .B2(new_n776_), .ZN(new_n818_));
  AOI211_X1 g617(.A(KEYINPUT114), .B(new_n775_), .C1(new_n600_), .C2(new_n608_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n808_), .A2(new_n607_), .B1(KEYINPUT112), .B2(KEYINPUT56), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n538_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n564_), .B1(new_n817_), .B2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n716_), .A2(new_n461_), .A3(new_n564_), .A4(new_n542_), .ZN(new_n826_));
  XOR2_X1   g625(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n826_), .B(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n248_), .B(new_n768_), .C1(new_n825_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n715_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n805_), .A2(new_n806_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n792_), .B1(new_n834_), .B2(new_n588_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n607_), .B1(new_n835_), .B2(new_n791_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n812_), .B1(new_n836_), .B2(new_n810_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n811_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n814_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n684_), .A3(new_n816_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n823_), .B2(KEYINPUT57), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n802_), .A2(new_n803_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n563_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n826_), .B(new_n827_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n249_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT115), .B1(new_n843_), .B2(new_n844_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n845_), .B(new_n768_), .C1(new_n846_), .C2(KEYINPUT59), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n825_), .B2(new_n829_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n830_), .A2(new_n848_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n461_), .B1(new_n847_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n833_), .B1(new_n852_), .B2(new_n832_), .ZN(G1340gat));
  NAND2_X1  g652(.A1(new_n847_), .A2(new_n851_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT116), .B(G120gat), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n716_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n716_), .B1(new_n831_), .B2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n831_), .A2(new_n855_), .A3(new_n858_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n854_), .A2(new_n859_), .B1(new_n860_), .B2(new_n856_), .ZN(G1341gat));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(G127gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n564_), .A2(KEYINPUT117), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(G127gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n854_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867_));
  AOI21_X1  g666(.A(G127gat), .B1(new_n831_), .B2(new_n564_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n865_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n847_), .B2(new_n851_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT118), .B1(new_n872_), .B2(new_n868_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(G1342gat));
  INV_X1    g673(.A(G134gat), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n542_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n854_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G134gat), .B1(new_n831_), .B2(new_n538_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(KEYINPUT119), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881_));
  INV_X1    g680(.A(new_n876_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n847_), .B2(new_n851_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n883_), .B2(new_n878_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n880_), .A2(new_n884_), .ZN(G1343gat));
  NOR3_X1   g684(.A1(new_n645_), .A2(new_n377_), .A3(new_n351_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n845_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n461_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n211_), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n716_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n212_), .ZN(G1345gat));
  AND2_X1   g690(.A1(new_n845_), .A2(new_n886_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n564_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT120), .B1(new_n887_), .B2(new_n563_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1346gat));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n207_), .A3(new_n538_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G162gat), .B1(new_n887_), .B2(new_n542_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1347gat));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  INV_X1    g702(.A(G169gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n375_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n292_), .A2(new_n380_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n715_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n904_), .B1(new_n905_), .B2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT62), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n905_), .A2(new_n259_), .A3(new_n908_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n909_), .B2(KEYINPUT62), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n903_), .B1(new_n911_), .B2(new_n913_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n909_), .A2(KEYINPUT62), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n915_), .A2(KEYINPUT121), .A3(new_n910_), .A4(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1348gat));
  AND2_X1   g716(.A1(new_n905_), .A2(new_n906_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n716_), .B1(KEYINPUT122), .B2(new_n260_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n260_), .A2(KEYINPUT122), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1349gat));
  AOI21_X1  g721(.A(new_n265_), .B1(new_n918_), .B2(new_n564_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n918_), .A2(new_n564_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n320_), .B2(new_n924_), .ZN(G1350gat));
  INV_X1    g724(.A(new_n278_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n918_), .A2(new_n926_), .A3(new_n538_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n918_), .A2(new_n684_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n928_), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(KEYINPUT123), .B1(new_n928_), .B2(G190gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n927_), .B1(new_n929_), .B2(new_n930_), .ZN(G1351gat));
  NAND3_X1  g730(.A1(new_n414_), .A2(new_n381_), .A3(new_n351_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n932_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n933_), .A2(G197gat), .A3(new_n715_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n933_), .A2(new_n715_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n303_), .ZN(new_n939_));
  AOI211_X1 g738(.A(KEYINPUT125), .B(G197gat), .C1(new_n933_), .C2(new_n715_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n936_), .A2(new_n939_), .A3(new_n940_), .ZN(G1352gat));
  NAND2_X1  g740(.A1(new_n933_), .A2(new_n613_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(G204gat), .ZN(new_n943_));
  INV_X1    g742(.A(new_n933_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n716_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n943_), .A2(KEYINPUT126), .B1(new_n945_), .B2(new_n302_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(KEYINPUT126), .B2(new_n943_), .ZN(G1353gat));
  NAND2_X1  g746(.A1(new_n933_), .A2(new_n564_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  AND2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n948_), .A2(new_n949_), .A3(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n948_), .B2(new_n949_), .ZN(G1354gat));
  AND3_X1   g751(.A1(new_n933_), .A2(G218gat), .A3(new_n684_), .ZN(new_n953_));
  AOI21_X1  g752(.A(KEYINPUT127), .B1(new_n933_), .B2(new_n538_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(G218gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n933_), .A2(KEYINPUT127), .A3(new_n538_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n953_), .B1(new_n955_), .B2(new_n956_), .ZN(G1355gat));
endmodule


