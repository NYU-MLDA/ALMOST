//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND4_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .A4(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT7), .ZN(new_n207_));
  OAI22_X1  g006(.A1(new_n207_), .A2(KEYINPUT64), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n203_), .A2(KEYINPUT7), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  AND3_X1   g009(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n215_), .A3(new_n221_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT65), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n224_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n220_), .B1(new_n230_), .B2(new_n210_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n222_), .B1(new_n231_), .B2(new_n215_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n205_), .A3(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n218_), .A2(KEYINPUT9), .A3(new_n219_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n213_), .A2(new_n235_), .A3(new_n236_), .A4(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G64gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT11), .Z(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT66), .B(G71gat), .ZN(new_n242_));
  INV_X1    g041(.A(G78gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT12), .B1(new_n239_), .B2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT67), .B(new_n222_), .C1(new_n231_), .C2(new_n215_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT65), .B1(new_n211_), .B2(new_n212_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n227_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n210_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n215_), .B1(new_n254_), .B2(new_n221_), .ZN(new_n255_));
  AOI211_X1 g054(.A(KEYINPUT8), .B(new_n220_), .C1(new_n210_), .C2(new_n213_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n251_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n238_), .B(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n250_), .A2(new_n257_), .A3(KEYINPUT69), .A4(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n248_), .A2(KEYINPUT12), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n249_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n239_), .B2(new_n248_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n202_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n265_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n272_));
  NOR4_X1   g071(.A1(new_n272_), .A2(KEYINPUT70), .A3(new_n249_), .A4(new_n269_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n239_), .A2(new_n248_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n239_), .A2(new_n248_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n268_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n271_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n278_), .A2(KEYINPUT72), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n238_), .B(KEYINPUT68), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n232_), .B2(new_n251_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n287_), .B2(new_n250_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n263_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n266_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n249_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n270_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT70), .ZN(new_n293_));
  INV_X1    g092(.A(new_n277_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n267_), .A2(new_n202_), .A3(new_n270_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n285_), .B1(new_n296_), .B2(new_n282_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .A4(new_n283_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n284_), .A2(new_n297_), .A3(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT72), .B1(new_n278_), .B2(new_n283_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n296_), .A2(new_n285_), .A3(new_n282_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n302_), .A2(new_n303_), .B1(new_n299_), .B2(new_n298_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT13), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n300_), .B1(new_n284_), .B2(new_n297_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n302_), .A2(new_n299_), .A3(new_n298_), .A4(new_n303_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT13), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313_));
  INV_X1    g112(.A(G1gat), .ZN(new_n314_));
  INV_X1    g113(.A(G8gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT14), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G1gat), .B(G8gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G43gat), .B(G50gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(G29gat), .B(G36gat), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n319_), .B(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n319_), .A2(new_n324_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n324_), .B(KEYINPUT15), .Z(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(new_n319_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G229gat), .A2(G233gat), .ZN(new_n329_));
  MUX2_X1   g128(.A(new_n325_), .B(new_n328_), .S(new_n329_), .Z(new_n330_));
  XNOR2_X1  g129(.A(G113gat), .B(G141gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G169gat), .B(G197gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT79), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n330_), .B(new_n335_), .Z(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT0), .ZN(new_n338_));
  INV_X1    g137(.A(G57gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(new_n216_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT90), .ZN(new_n343_));
  OAI22_X1  g142(.A1(new_n343_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(KEYINPUT90), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT2), .ZN(new_n348_));
  INV_X1    g147(.A(G141gat), .ZN(new_n349_));
  INV_X1    g148(.A(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n343_), .A3(KEYINPUT3), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n346_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT89), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n354_), .B(KEYINPUT89), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n356_), .B(KEYINPUT1), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n347_), .B(new_n351_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G127gat), .B(G134gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G113gat), .B(G120gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(KEYINPUT4), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n364_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(KEYINPUT4), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT101), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n369_), .ZN(new_n371_));
  AOI211_X1 g170(.A(new_n342_), .B(new_n366_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n365_), .A2(new_n367_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n342_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n341_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n370_), .A2(new_n371_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n366_), .A2(new_n342_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n375_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n341_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n376_), .B1(new_n381_), .B2(KEYINPUT102), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(KEYINPUT102), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(G183gat), .A3(G190gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G183gat), .ZN(new_n389_));
  INV_X1    g188(.A(G190gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT23), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n387_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT80), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT24), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT26), .B(G190gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT25), .B(G183gat), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n395_), .A2(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n394_), .B(KEYINPUT80), .Z(new_n400_));
  NAND2_X1  g199(.A1(G169gat), .A2(G176gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n393_), .B(new_n399_), .C1(new_n402_), .C2(new_n396_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n391_), .A2(new_n386_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(G183gat), .B2(G190gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n401_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT22), .B(G169gat), .ZN(new_n407_));
  INV_X1    g206(.A(G176gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT82), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n403_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n411_), .B(KEYINPUT83), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT30), .ZN(new_n417_));
  XOR2_X1   g216(.A(G15gat), .B(G43gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT84), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G227gat), .A2(G233gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n422_), .B(KEYINPUT85), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n421_), .B(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n415_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT88), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n415_), .A2(new_n417_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n424_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n415_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n364_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n364_), .A2(new_n434_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n435_), .A2(new_n436_), .A3(KEYINPUT86), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n427_), .A2(new_n433_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n427_), .B2(new_n433_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n361_), .A2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n442_), .B(KEYINPUT28), .Z(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G228gat), .A2(G233gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT92), .B(G204gat), .Z(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G197gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT91), .B(G197gat), .Z(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G204gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT94), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT21), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G211gat), .B(G218gat), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n449_), .A2(G204gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n447_), .A2(G197gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT21), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT93), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n448_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n461_), .A2(new_n454_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n361_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n446_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n446_), .B1(new_n361_), .B2(new_n441_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n455_), .B2(new_n463_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n445_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n470_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n445_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n455_), .A2(new_n463_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n472_), .B(new_n473_), .C1(new_n446_), .C2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G22gat), .B(G50gat), .Z(new_n476_));
  AND3_X1   g275(.A1(new_n471_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n444_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n475_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n476_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n471_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n443_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n440_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n479_), .B(new_n484_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n384_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n401_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n407_), .B(KEYINPUT98), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(new_n408_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n393_), .B1(G183gat), .B2(G190gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT99), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n491_), .A2(KEYINPUT99), .A3(new_n492_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n398_), .B(KEYINPUT96), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n397_), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n499_));
  AOI22_X1  g298(.A1(new_n499_), .A2(new_n394_), .B1(new_n386_), .B2(new_n391_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n498_), .B(new_n500_), .C1(new_n402_), .C2(new_n499_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n495_), .A2(new_n496_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n464_), .A2(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n503_), .B(KEYINPUT20), .C1(new_n464_), .C2(new_n413_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G226gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT19), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n413_), .A2(new_n464_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n508_), .B(new_n510_), .C1(new_n464_), .C2(new_n502_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G8gat), .B(G36gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT18), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G64gat), .B(G92gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  NAND3_X1  g314(.A1(new_n507_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n516_), .B1(new_n517_), .B2(KEYINPUT100), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n507_), .A2(new_n511_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT100), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n515_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT27), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n515_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n504_), .A2(new_n506_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n506_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n464_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n501_), .A2(new_n493_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n509_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n525_), .B1(new_n528_), .B2(new_n508_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n523_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n530_), .A2(KEYINPUT27), .A3(new_n516_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n522_), .A2(new_n531_), .ZN(new_n532_));
  AOI211_X1 g331(.A(new_n375_), .B(new_n341_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n533_), .A2(KEYINPUT33), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n341_), .B1(new_n373_), .B2(new_n342_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n366_), .A2(new_n374_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n377_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n533_), .B2(KEYINPUT33), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n518_), .A2(new_n534_), .A3(new_n521_), .A4(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n382_), .A2(new_n383_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n519_), .B1(new_n541_), .B2(new_n523_), .ZN(new_n542_));
  OAI211_X1 g341(.A(KEYINPUT32), .B(new_n515_), .C1(new_n524_), .C2(new_n529_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n539_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n485_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(new_n440_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n488_), .A2(new_n532_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n239_), .A2(new_n324_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT34), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT35), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n549_), .A2(KEYINPUT75), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n264_), .A2(new_n327_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n552_), .A2(new_n553_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n556_), .B(new_n555_), .C1(new_n553_), .C2(new_n552_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT74), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT36), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n565_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n559_), .A2(new_n569_), .A3(new_n560_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n570_), .B2(KEYINPUT76), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n567_), .B(new_n570_), .C1(KEYINPUT76), .C2(new_n572_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT16), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT17), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT77), .Z(new_n582_));
  INV_X1    g381(.A(new_n248_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n319_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n583_), .B(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n582_), .A2(KEYINPUT78), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n580_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT17), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT78), .B1(new_n582_), .B2(new_n586_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n576_), .A2(new_n592_), .ZN(new_n593_));
  NOR4_X1   g392(.A1(new_n312_), .A2(new_n336_), .A3(new_n548_), .A4(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n314_), .A3(new_n384_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT38), .Z(new_n596_));
  INV_X1    g395(.A(new_n310_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(new_n336_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n548_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n592_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n571_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n314_), .B1(new_n604_), .B2(new_n384_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n596_), .A2(new_n605_), .ZN(G1324gat));
  XNOR2_X1  g405(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n607_));
  INV_X1    g406(.A(new_n532_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n603_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(G8gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT39), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n594_), .A2(new_n315_), .A3(new_n608_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n607_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(KEYINPUT39), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n609_), .B2(G8gat), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n612_), .B(new_n607_), .C1(new_n614_), .C2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n613_), .A2(new_n618_), .ZN(G1325gat));
  NAND2_X1  g418(.A1(new_n604_), .A2(new_n440_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G15gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT41), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT41), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n623_), .A3(G15gat), .ZN(new_n624_));
  INV_X1    g423(.A(G15gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n594_), .A2(new_n625_), .A3(new_n440_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT104), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n622_), .A2(new_n629_), .A3(new_n624_), .A4(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(G1326gat));
  XOR2_X1   g430(.A(new_n485_), .B(KEYINPUT105), .Z(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(G22gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT106), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n594_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n604_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G22gat), .B1(new_n637_), .B2(new_n633_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(KEYINPUT42), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(KEYINPUT42), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(G1327gat));
  NOR2_X1   g440(.A1(new_n592_), .A2(new_n571_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n600_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G29gat), .B1(new_n644_), .B2(new_n384_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n647_), .B(KEYINPUT43), .C1(new_n548_), .C2(new_n576_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n486_), .A2(new_n487_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n532_), .A3(new_n540_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n545_), .A2(new_n547_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  INV_X1    g452(.A(new_n576_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n654_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n647_), .B1(new_n657_), .B2(KEYINPUT43), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n599_), .A2(new_n592_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n646_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n662_), .A2(G29gat), .A3(new_n384_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n660_), .B(KEYINPUT44), .C1(new_n656_), .C2(new_n658_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n645_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n662_), .A2(new_n608_), .A3(new_n664_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n600_), .A2(new_n668_), .A3(new_n608_), .A4(new_n642_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n667_), .B1(new_n672_), .B2(KEYINPUT45), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n673_), .B1(KEYINPUT45), .B2(new_n672_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n670_), .A2(new_n671_), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n670_), .B2(new_n674_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  NAND4_X1  g476(.A1(new_n662_), .A2(G43gat), .A3(new_n440_), .A4(new_n664_), .ZN(new_n678_));
  INV_X1    g477(.A(G43gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n440_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n643_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g482(.A(G50gat), .B1(new_n644_), .B2(new_n632_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n662_), .A2(G50gat), .A3(new_n546_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n664_), .ZN(G1331gat));
  INV_X1    g485(.A(new_n336_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n548_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n593_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n597_), .A2(KEYINPUT110), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT110), .B1(new_n597_), .B2(new_n689_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n339_), .B1(new_n695_), .B2(new_n540_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n312_), .A2(new_n688_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n697_), .A2(G57gat), .A3(new_n384_), .A4(new_n603_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT112), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n696_), .A2(KEYINPUT112), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1332gat));
  NAND2_X1  g502(.A1(new_n697_), .A2(new_n603_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G64gat), .B1(new_n704_), .B2(new_n532_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT48), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n532_), .A2(G64gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n695_), .B2(new_n707_), .ZN(G1333gat));
  OAI21_X1  g507(.A(G71gat), .B1(new_n704_), .B2(new_n680_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT49), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n680_), .A2(G71gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n695_), .B2(new_n711_), .ZN(G1334gat));
  OAI21_X1  g511(.A(G78gat), .B1(new_n704_), .B2(new_n633_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT50), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n632_), .A2(new_n243_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n695_), .B2(new_n715_), .ZN(G1335gat));
  NOR3_X1   g515(.A1(new_n310_), .A2(new_n592_), .A3(new_n687_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n540_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n312_), .A2(new_n642_), .A3(new_n688_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT113), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n384_), .A2(new_n216_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(G1336gat));
  OAI21_X1  g522(.A(G92gat), .B1(new_n718_), .B2(new_n532_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n608_), .A2(new_n217_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n721_), .B2(new_n725_), .ZN(G1337gat));
  OAI211_X1 g525(.A(new_n440_), .B(new_n717_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G99gat), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n440_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n697_), .A2(KEYINPUT113), .A3(new_n642_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n720_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n730_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT115), .B1(new_n729_), .B2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT115), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n728_), .B(new_n737_), .C1(new_n721_), .C2(new_n730_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n735_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n736_), .B1(new_n735_), .B2(new_n738_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1338gat));
  OAI21_X1  g540(.A(G106gat), .B1(new_n718_), .B2(new_n485_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n546_), .A2(new_n205_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n721_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT53), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n742_), .A2(KEYINPUT52), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n742_), .A2(KEYINPUT52), .ZN(new_n750_));
  OAI221_X1 g549(.A(new_n748_), .B1(new_n721_), .B2(new_n745_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n747_), .A2(new_n751_), .ZN(G1339gat));
  NOR2_X1   g551(.A1(new_n608_), .A2(new_n540_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n486_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n293_), .A2(new_n757_), .A3(new_n295_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n267_), .A2(new_n275_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n268_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n272_), .A2(new_n249_), .A3(new_n269_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n759_), .A2(new_n760_), .B1(new_n761_), .B2(KEYINPUT55), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(KEYINPUT56), .A4(new_n282_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n298_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n336_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n763_), .B2(new_n282_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n769_), .A2(new_n764_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n763_), .A2(KEYINPUT56), .A3(new_n282_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n330_), .A2(new_n334_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n328_), .A2(G229gat), .A3(G233gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n325_), .A2(new_n329_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n334_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT57), .B(new_n571_), .C1(new_n772_), .C2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT117), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n271_), .A2(new_n273_), .A3(KEYINPUT55), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n272_), .A2(new_n274_), .A3(new_n249_), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n757_), .A2(new_n292_), .B1(new_n782_), .B2(new_n268_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n282_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(KEYINPUT116), .A3(new_n771_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n777_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n602_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(KEYINPUT57), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n780_), .A2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n766_), .A2(new_n777_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n785_), .B(new_n283_), .C1(new_n758_), .C2(new_n762_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT58), .B(new_n795_), .C1(new_n769_), .C2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n654_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n786_), .A2(new_n771_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT58), .B1(new_n799_), .B2(new_n795_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n571_), .B1(new_n772_), .B2(new_n778_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n592_), .B1(new_n794_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n593_), .A2(new_n687_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n310_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n687_), .B(new_n756_), .C1(new_n805_), .C2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(KEYINPUT118), .A3(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n687_), .A2(G113gat), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n779_), .A2(KEYINPUT117), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n792_), .B1(new_n791_), .B2(KEYINPUT57), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n804_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n809_), .B1(new_n821_), .B2(new_n601_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n822_), .B2(new_n755_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT59), .B(new_n756_), .C1(new_n805_), .C2(new_n809_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n817_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT119), .B1(new_n816_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n825_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n815_), .A4(new_n814_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(G1340gat));
  NOR2_X1   g629(.A1(new_n822_), .A2(new_n755_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n832_));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n597_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT120), .ZN(new_n837_));
  INV_X1    g636(.A(new_n312_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n833_), .B2(new_n839_), .ZN(G1341gat));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n831_), .A2(new_n841_), .A3(new_n592_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n601_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n841_), .ZN(G1342gat));
  INV_X1    g643(.A(G134gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n831_), .A2(new_n845_), .A3(new_n602_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n576_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n845_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n846_), .B(KEYINPUT121), .C1(new_n847_), .C2(new_n845_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1343gat));
  NAND2_X1  g651(.A1(new_n821_), .A2(new_n601_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n809_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n487_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n753_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n336_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n349_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n838_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n350_), .ZN(G1345gat));
  OAI21_X1  g660(.A(KEYINPUT122), .B1(new_n857_), .B2(new_n601_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n822_), .A2(new_n487_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n592_), .A4(new_n753_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n862_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n857_), .B2(new_n576_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n571_), .A2(G162gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n857_), .B2(new_n871_), .ZN(G1347gat));
  NOR4_X1   g671(.A1(new_n632_), .A2(new_n384_), .A3(new_n532_), .A4(new_n680_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n855_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT124), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n855_), .A2(new_n876_), .A3(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n687_), .A3(new_n490_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n855_), .A2(new_n687_), .A3(new_n873_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n881_), .A3(G169gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n880_), .B2(G169gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(KEYINPUT123), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885_));
  AOI211_X1 g684(.A(new_n885_), .B(new_n881_), .C1(new_n880_), .C2(G169gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n879_), .B1(new_n884_), .B2(new_n886_), .ZN(G1348gat));
  NAND2_X1  g686(.A1(new_n878_), .A2(new_n597_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n822_), .A2(new_n384_), .A3(new_n532_), .A4(new_n486_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n838_), .A2(new_n408_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n889_), .A2(KEYINPUT125), .A3(new_n890_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n888_), .A2(new_n408_), .B1(new_n893_), .B2(new_n894_), .ZN(G1349gat));
  AOI21_X1  g694(.A(G183gat), .B1(new_n889_), .B2(new_n592_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n601_), .A2(new_n497_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n878_), .B2(new_n897_), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n878_), .A2(new_n602_), .A3(new_n397_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n576_), .B1(new_n875_), .B2(new_n877_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n390_), .B2(new_n900_), .ZN(G1351gat));
  NOR2_X1   g700(.A1(new_n532_), .A2(new_n384_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n863_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n336_), .ZN(new_n904_));
  INV_X1    g703(.A(G197gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1352gat));
  NAND3_X1  g705(.A1(new_n863_), .A2(new_n312_), .A3(new_n902_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n447_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT126), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n907_), .B2(G204gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n909_), .B2(new_n912_), .ZN(G1353gat));
  NOR2_X1   g712(.A1(new_n903_), .A2(new_n601_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  AND2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n914_), .B2(new_n915_), .ZN(G1354gat));
  INV_X1    g717(.A(new_n903_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G218gat), .B1(new_n919_), .B2(new_n602_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n654_), .A2(G218gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n919_), .B2(new_n922_), .ZN(G1355gat));
endmodule


