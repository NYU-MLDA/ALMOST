//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(new_n207_), .A3(KEYINPUT87), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(KEYINPUT3), .B2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(KEYINPUT3), .B2(new_n208_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G155gat), .B(G162gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n206_), .A2(new_n207_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n203_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT86), .ZN(new_n222_));
  XOR2_X1   g021(.A(G113gat), .B(G120gat), .Z(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n218_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n224_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(KEYINPUT4), .A3(new_n228_), .ZN(new_n229_));
  OR3_X1    g028(.A1(new_n227_), .A2(new_n224_), .A3(KEYINPUT4), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n202_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G1gat), .B(G29gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G85gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT0), .B(G57gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  INV_X1    g034(.A(new_n202_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n231_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n235_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G226gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT19), .ZN(new_n242_));
  INV_X1    g041(.A(G183gat), .ZN(new_n243_));
  INV_X1    g042(.A(G190gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT23), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT23), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G183gat), .A3(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT81), .Z(new_n252_));
  OR2_X1    g051(.A1(new_n252_), .A2(KEYINPUT24), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT80), .B1(new_n243_), .B2(KEYINPUT25), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT25), .B(G183gat), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n254_), .B(new_n255_), .C1(new_n256_), .C2(KEYINPUT80), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n252_), .A2(KEYINPUT24), .A3(new_n258_), .ZN(new_n259_));
  AND4_X1   g058(.A1(new_n250_), .A2(new_n253_), .A3(new_n257_), .A4(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT22), .B(G169gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(KEYINPUT83), .ZN(new_n262_));
  INV_X1    g061(.A(G169gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT83), .B1(new_n263_), .B2(KEYINPUT22), .ZN(new_n264_));
  INV_X1    g063(.A(G176gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n258_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(KEYINPUT84), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n245_), .A2(new_n249_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n243_), .A2(new_n244_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT85), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n267_), .A2(KEYINPUT84), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n260_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G197gat), .B(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(KEYINPUT90), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(KEYINPUT90), .A3(new_n278_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n277_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n280_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n281_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n275_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n250_), .A2(new_n270_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n261_), .A2(new_n265_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n258_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n256_), .A2(new_n255_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT24), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n251_), .A2(new_n294_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n259_), .A2(new_n269_), .A3(new_n293_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT20), .B1(new_n297_), .B2(new_n287_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n242_), .B1(new_n289_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT20), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n275_), .B2(new_n288_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT94), .B1(new_n297_), .B2(new_n287_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n297_), .A2(KEYINPUT94), .A3(new_n287_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n299_), .B1(new_n305_), .B2(new_n242_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G8gat), .B(G36gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT18), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G64gat), .B(G92gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n308_), .B(new_n309_), .Z(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT32), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n305_), .A2(new_n242_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n289_), .A2(new_n242_), .A3(new_n298_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n316_), .A3(new_n311_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n240_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n310_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n242_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n304_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(new_n302_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n322_), .B2(new_n301_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n319_), .B1(new_n323_), .B2(new_n315_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n314_), .A2(new_n316_), .A3(new_n310_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT95), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n314_), .A2(new_n316_), .A3(KEYINPUT95), .A4(new_n310_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT33), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n239_), .A2(KEYINPUT96), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n226_), .A2(new_n228_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT97), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT97), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n226_), .A2(new_n334_), .A3(new_n228_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n236_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n229_), .A2(new_n202_), .A3(new_n230_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n235_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n239_), .B2(new_n330_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT96), .B1(new_n239_), .B2(new_n330_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n331_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n318_), .B1(new_n329_), .B2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G22gat), .B(G50gat), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n220_), .A2(KEYINPUT29), .ZN(new_n346_));
  XOR2_X1   g145(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n220_), .A2(KEYINPUT29), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n345_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n347_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n350_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n344_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT89), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n352_), .A2(KEYINPUT89), .A3(new_n355_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n288_), .B1(new_n220_), .B2(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G228gat), .A2(G233gat), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n361_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364_));
  OR3_X1    g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(KEYINPUT92), .B(new_n364_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n360_), .B(new_n361_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT92), .B1(new_n368_), .B2(new_n364_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n358_), .B(new_n359_), .C1(new_n367_), .C2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n364_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT93), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT93), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n368_), .A2(new_n373_), .A3(new_n364_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n372_), .A2(new_n374_), .A3(new_n356_), .A4(new_n365_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n327_), .A2(new_n377_), .A3(new_n328_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n306_), .A2(new_n319_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n325_), .A3(KEYINPUT27), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n240_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n382_), .ZN(new_n383_));
  OAI22_X1  g182(.A1(new_n343_), .A2(new_n376_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385_));
  INV_X1    g184(.A(G43gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n275_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n275_), .A2(new_n388_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n224_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n224_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(G15gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT31), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n396_), .A2(new_n401_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n381_), .A2(new_n376_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n240_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n384_), .A2(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G85gat), .B(G92gat), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(KEYINPUT8), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT7), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n411_), .B(new_n412_), .C1(G99gat), .C2(G106gat), .ZN(new_n413_));
  INV_X1    g212(.A(G99gat), .ZN(new_n414_));
  INV_X1    g213(.A(G106gat), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n414_), .B(new_n415_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G99gat), .A2(G106gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT6), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(G99gat), .A3(G106gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n410_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(KEYINPUT66), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT66), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n413_), .A2(new_n416_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n427_), .A3(new_n422_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(KEYINPUT67), .A3(new_n408_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT8), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT67), .B1(new_n428_), .B2(new_n408_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n424_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT10), .B(G99gat), .Z(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n415_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n408_), .A2(KEYINPUT9), .ZN(new_n435_));
  INV_X1    g234(.A(G85gat), .ZN(new_n436_));
  INV_X1    g235(.A(G92gat), .ZN(new_n437_));
  OR3_X1    g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT9), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n434_), .A2(new_n435_), .A3(new_n422_), .A4(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G57gat), .B(G64gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G71gat), .B(G78gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT11), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n440_), .A2(KEYINPUT11), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n443_), .A2(new_n441_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n440_), .A2(KEYINPUT11), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n442_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n432_), .A2(new_n439_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT68), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n432_), .A2(new_n439_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n432_), .A2(new_n452_), .A3(new_n439_), .A4(new_n446_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n448_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G230gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT64), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n439_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT8), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n417_), .A2(KEYINPUT66), .B1(new_n419_), .B2(new_n421_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n409_), .B1(new_n460_), .B2(new_n427_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n461_), .B2(KEYINPUT67), .ZN(new_n462_));
  INV_X1    g261(.A(new_n431_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n458_), .B1(new_n464_), .B2(new_n424_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n456_), .B1(new_n465_), .B2(new_n446_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT12), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n468_));
  AOI211_X1 g267(.A(KEYINPUT12), .B(new_n446_), .C1(new_n432_), .C2(new_n439_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n466_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n457_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G120gat), .B(G148gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(G176gat), .B(G204gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT70), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n457_), .A2(new_n470_), .A3(new_n476_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(KEYINPUT70), .A3(new_n477_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT13), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(KEYINPUT13), .A3(new_n482_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G1gat), .ZN(new_n487_));
  INV_X1    g286(.A(G8gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT74), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(KEYINPUT74), .B(KEYINPUT14), .C1(new_n487_), .C2(new_n488_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G1gat), .B(G8gat), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n491_), .A2(new_n495_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G29gat), .B(G36gat), .Z(new_n501_));
  XOR2_X1   g300(.A(G43gat), .B(G50gat), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(KEYINPUT75), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n506_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT75), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n500_), .A2(KEYINPUT76), .A3(new_n507_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n507_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n512_), .B1(new_n513_), .B2(new_n499_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n508_), .B(KEYINPUT15), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(new_n499_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(KEYINPUT78), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n499_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT77), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n513_), .A2(KEYINPUT77), .A3(new_n499_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n523_), .A2(new_n524_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n525_), .B2(new_n516_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT78), .B1(new_n515_), .B2(new_n519_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT79), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G169gat), .B(G197gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(KEYINPUT79), .B(new_n531_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n486_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n407_), .A2(new_n536_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n462_), .A2(new_n463_), .B1(new_n423_), .B2(new_n410_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n518_), .B1(new_n538_), .B2(new_n458_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n432_), .A2(new_n439_), .A3(new_n508_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(KEYINPUT71), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n432_), .A2(new_n439_), .A3(new_n508_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n518_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n432_), .B2(new_n439_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n547_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n539_), .A2(KEYINPUT71), .A3(new_n540_), .A4(new_n544_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT72), .B1(new_n546_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT36), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n541_), .A2(new_n545_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT72), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n554_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n553_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n567_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n564_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n567_), .B2(new_n559_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT37), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT73), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n446_), .B(new_n499_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT16), .ZN(new_n582_));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n579_), .A2(new_n580_), .A3(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(KEYINPUT17), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n579_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n576_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n537_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n487_), .A3(new_n240_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT98), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n590_), .A2(new_n593_), .A3(new_n487_), .A4(new_n240_), .ZN(new_n594_));
  XOR2_X1   g393(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT100), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n562_), .A2(new_n565_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT102), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n407_), .A2(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n481_), .A2(KEYINPUT13), .A3(new_n482_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n483_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n535_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT101), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n536_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n602_), .A2(new_n587_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n487_), .B1(new_n612_), .B2(new_n240_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n592_), .A2(new_n594_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n614_), .B2(new_n595_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n598_), .A2(new_n615_), .ZN(G1324gat));
  NAND3_X1  g415(.A1(new_n590_), .A2(new_n488_), .A3(new_n381_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT103), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n381_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n620_));
  AND4_X1   g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .A4(G8gat), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n488_), .B1(KEYINPUT103), .B2(KEYINPUT39), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n619_), .A2(new_n622_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n617_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT40), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT40), .B(new_n617_), .C1(new_n621_), .C2(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(G1325gat));
  INV_X1    g427(.A(new_n404_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n612_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT104), .B1(new_n631_), .B2(new_n398_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n633_), .A3(G15gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n632_), .A2(KEYINPUT41), .A3(new_n634_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n590_), .A2(new_n398_), .A3(new_n629_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(G1326gat));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n590_), .A2(new_n641_), .A3(new_n376_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT42), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n612_), .A2(new_n376_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(G22gat), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT42), .B(new_n641_), .C1(new_n612_), .C2(new_n376_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(new_n599_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n588_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT106), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n537_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n240_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n606_), .A2(KEYINPUT101), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n536_), .A2(new_n608_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n588_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n384_), .A2(new_n404_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n405_), .A2(new_n406_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n576_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n573_), .A2(new_n575_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n407_), .B2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n656_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n587_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n660_), .B1(new_n659_), .B2(new_n576_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n407_), .A2(KEYINPUT43), .A3(new_n662_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n667_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n666_), .A2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n240_), .A2(G29gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n653_), .B1(new_n671_), .B2(new_n672_), .ZN(G1328gat));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n670_), .B(new_n381_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G36gat), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n537_), .A2(new_n680_), .A3(new_n381_), .A4(new_n650_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n676_), .B(new_n677_), .C1(new_n679_), .C2(new_n683_), .ZN(new_n684_));
  AND4_X1   g483(.A1(new_n674_), .A2(new_n679_), .A3(new_n675_), .A4(new_n683_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1329gat));
  NOR2_X1   g485(.A1(new_n404_), .A2(new_n386_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n666_), .A2(KEYINPUT109), .A3(new_n670_), .A4(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT110), .B(G43gat), .Z(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n651_), .B2(new_n404_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n670_), .B(new_n687_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n688_), .A2(new_n692_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT47), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n688_), .A2(new_n692_), .A3(new_n695_), .A4(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1330gat));
  AOI211_X1 g499(.A(G50gat), .B(new_n651_), .C1(new_n375_), .C2(new_n370_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n670_), .B(new_n376_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(G50gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT112), .ZN(G1331gat));
  NAND2_X1  g503(.A1(new_n589_), .A2(new_n604_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(KEYINPUT113), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n407_), .A2(new_n535_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(KEYINPUT113), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(G57gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n240_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n588_), .A2(new_n535_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n486_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n602_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n382_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n712_), .A2(new_n718_), .ZN(G1332gat));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n716_), .B2(new_n381_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT48), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n710_), .A2(new_n720_), .A3(new_n381_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1333gat));
  INV_X1    g523(.A(G71gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n716_), .B2(new_n629_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT49), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n710_), .A2(new_n725_), .A3(new_n629_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n716_), .B2(new_n376_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT114), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n731_), .A2(new_n732_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735_));
  OR3_X1    g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n710_), .A2(new_n730_), .A3(new_n376_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(G1335gat));
  NAND2_X1  g538(.A1(new_n661_), .A2(new_n663_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n486_), .A2(new_n587_), .A3(new_n535_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742_), .B2(new_n382_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n708_), .A2(new_n604_), .A3(new_n650_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n436_), .A3(new_n240_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1336gat));
  NAND3_X1  g545(.A1(new_n744_), .A2(new_n437_), .A3(new_n381_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n437_), .ZN(G1337gat));
  NAND3_X1  g548(.A1(new_n744_), .A2(new_n433_), .A3(new_n629_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n742_), .A2(new_n404_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n414_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(KEYINPUT115), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n752_), .B(new_n754_), .ZN(G1338gat));
  NAND3_X1  g554(.A1(new_n744_), .A2(new_n415_), .A3(new_n376_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n740_), .A2(new_n376_), .A3(new_n741_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(G106gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G106gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g561(.A(KEYINPUT121), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT59), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT58), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n468_), .A2(new_n469_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n448_), .A2(new_n453_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n456_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n470_), .A2(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n466_), .B(KEYINPUT55), .C1(new_n468_), .C2(new_n469_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n477_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n772_), .B2(new_n477_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(KEYINPUT118), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n477_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(KEYINPUT118), .A3(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n526_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n532_), .B1(new_n525_), .B2(new_n517_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(KEYINPUT117), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n516_), .B1(new_n518_), .B2(new_n499_), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n780_), .A2(KEYINPUT117), .B1(new_n515_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n779_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(new_n480_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n778_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n765_), .B1(new_n775_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n776_), .A2(new_n777_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n477_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT58), .A3(new_n778_), .A4(new_n785_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n576_), .A2(new_n787_), .A3(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n481_), .A2(new_n482_), .A3(new_n784_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n480_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n796_), .B2(KEYINPUT116), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(new_n795_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n648_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n793_), .B1(new_n800_), .B2(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n802_), .B(new_n648_), .C1(new_n797_), .C2(new_n799_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n588_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n713_), .B1(new_n603_), .B2(new_n483_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n662_), .B2(new_n807_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n576_), .A2(new_n806_), .A3(KEYINPUT54), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n804_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n404_), .A2(new_n382_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n405_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n764_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n814_), .A2(KEYINPUT120), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(KEYINPUT120), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n764_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n804_), .B2(new_n811_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n763_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n481_), .A2(new_n482_), .A3(new_n784_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n535_), .A2(new_n480_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n824_), .B2(new_n798_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n799_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n599_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n802_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n793_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n810_), .B1(new_n830_), .B2(new_n588_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT59), .B1(new_n831_), .B2(new_n814_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n820_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(KEYINPUT121), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n821_), .A2(new_n535_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G113gat), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n831_), .B2(new_n814_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n812_), .A2(KEYINPUT119), .A3(new_n815_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(G113gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n535_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n836_), .A2(new_n842_), .ZN(G1340gat));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n486_), .B2(KEYINPUT60), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(KEYINPUT60), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(KEYINPUT122), .B2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n840_), .B(new_n847_), .C1(KEYINPUT122), .C2(new_n845_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n816_), .A2(new_n486_), .A3(new_n820_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n844_), .ZN(G1341gat));
  NAND3_X1  g649(.A1(new_n838_), .A2(new_n839_), .A3(new_n587_), .ZN(new_n851_));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT123), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n855_), .A3(new_n852_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n816_), .A2(new_n763_), .A3(new_n820_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT121), .B1(new_n832_), .B2(new_n833_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n588_), .A2(new_n852_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n854_), .A2(new_n856_), .B1(new_n859_), .B2(new_n860_), .ZN(G1342gat));
  NAND3_X1  g660(.A1(new_n821_), .A2(new_n576_), .A3(new_n834_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G134gat), .ZN(new_n863_));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n840_), .A2(new_n864_), .A3(new_n601_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1343gat));
  NAND3_X1  g665(.A1(new_n404_), .A2(new_n376_), .A3(new_n240_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n831_), .A2(new_n381_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n535_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n604_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n587_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n868_), .A2(new_n876_), .A3(new_n601_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n868_), .B2(new_n576_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT124), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n868_), .A2(new_n576_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n881_), .B(new_n877_), .C1(new_n882_), .C2(new_n876_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(G1347gat));
  AND2_X1   g683(.A1(new_n812_), .A2(new_n381_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n404_), .A2(new_n376_), .A3(new_n240_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887_), .B2(new_n605_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n887_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n535_), .A3(new_n261_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT62), .B(G169gat), .C1(new_n887_), .C2(new_n605_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n892_), .A3(new_n893_), .ZN(G1348gat));
  NOR2_X1   g693(.A1(new_n887_), .A2(new_n486_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n265_), .ZN(G1349gat));
  NAND3_X1  g695(.A1(new_n885_), .A2(new_n587_), .A3(new_n886_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n256_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n243_), .B2(new_n897_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n887_), .B2(new_n662_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n601_), .A2(new_n255_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n887_), .B2(new_n901_), .ZN(G1351gat));
  NOR2_X1   g701(.A1(new_n629_), .A2(new_n383_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n885_), .A2(new_n535_), .A3(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g704(.A1(new_n885_), .A2(new_n903_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT125), .B(G204gat), .Z(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(new_n604_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n885_), .A2(new_n903_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n909_), .A2(new_n486_), .B1(new_n910_), .B2(G204gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n908_), .A2(new_n911_), .ZN(G1353gat));
  NAND4_X1  g711(.A1(new_n812_), .A2(new_n587_), .A3(new_n381_), .A4(new_n903_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT63), .B(G211gat), .Z(new_n914_));
  OR2_X1    g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n913_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1354gat));
  AOI21_X1  g719(.A(G218gat), .B1(new_n906_), .B2(new_n601_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n576_), .A2(G218gat), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT127), .Z(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n906_), .B2(new_n923_), .ZN(G1355gat));
endmodule


