//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n206_), .B(KEYINPUT71), .ZN(new_n211_));
  INV_X1    g010(.A(new_n209_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G29gat), .B(G36gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n214_), .B(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n218_), .A2(KEYINPUT72), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G229gat), .A2(G233gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(KEYINPUT72), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n217_), .B(KEYINPUT15), .Z(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n214_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n217_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n226_), .B(new_n220_), .C1(new_n214_), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G141gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G169gat), .B(G197gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n230_), .B(new_n231_), .Z(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n223_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G141gat), .A2(G148gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(KEYINPUT1), .B2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n242_), .A2(KEYINPUT1), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n240_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n238_), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n247_), .B1(new_n237_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n239_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n237_), .A2(new_n248_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n250_), .A2(new_n252_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n242_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(new_n241_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n245_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT28), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G22gat), .B(G50gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n261_), .A2(new_n263_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT80), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(G197gat), .B(G204gat), .Z(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(KEYINPUT81), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(G197gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT21), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  OAI221_X1 g076(.A(new_n271_), .B1(KEYINPUT21), .B2(new_n272_), .C1(new_n273_), .C2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n271_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(KEYINPUT21), .A3(new_n272_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n282_));
  AND2_X1   g081(.A1(G228gat), .A2(G233gat), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G78gat), .B(G106gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT82), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  OR3_X1    g087(.A1(new_n284_), .A2(new_n285_), .A3(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n267_), .A2(new_n270_), .A3(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n290_), .A2(KEYINPUT83), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n265_), .A2(new_n266_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(KEYINPUT83), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .A4(new_n289_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT20), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  MUX2_X1   g102(.A(new_n301_), .B(new_n303_), .S(KEYINPUT24), .Z(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n305_));
  INV_X1    g104(.A(G183gat), .ZN(new_n306_));
  INV_X1    g105(.A(G190gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT25), .B(G183gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT26), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(G190gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n313_), .B(new_n316_), .C1(new_n317_), .C2(new_n314_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n304_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n308_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n310_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n305_), .B2(new_n322_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n321_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n299_), .B1(new_n327_), .B2(new_n281_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n300_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n303_), .B2(new_n334_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n324_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n313_), .B(KEYINPUT86), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n338_), .A2(new_n317_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n325_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(G169gat), .ZN(new_n344_));
  INV_X1    g143(.A(G169gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n345_), .A2(KEYINPUT22), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT89), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(KEYINPUT22), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(G169gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT89), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(G176gat), .B1(new_n347_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n302_), .B(KEYINPUT88), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n352_), .A2(KEYINPUT90), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT90), .ZN(new_n355_));
  INV_X1    g154(.A(G176gat), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n350_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n353_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n355_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n342_), .B1(new_n354_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT91), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT90), .B1(new_n352_), .B2(new_n353_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT91), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n342_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n340_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n281_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n333_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT92), .B1(new_n369_), .B2(new_n370_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n340_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n367_), .B1(new_n366_), .B2(new_n342_), .ZN(new_n374_));
  AOI211_X1 g173(.A(KEYINPUT91), .B(new_n341_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n281_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n327_), .A2(new_n281_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT20), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n372_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n331_), .B(KEYINPUT85), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n371_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n385_), .A2(new_n390_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n298_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n298_), .B1(new_n385_), .B2(new_n390_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n373_), .A2(new_n370_), .A3(new_n362_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n332_), .B1(new_n395_), .B2(new_n328_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n372_), .A2(new_n378_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n397_), .B2(KEYINPUT96), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n376_), .A2(new_n281_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n380_), .B1(new_n399_), .B2(KEYINPUT92), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n378_), .A4(new_n383_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n390_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n394_), .B1(new_n403_), .B2(KEYINPUT97), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT97), .ZN(new_n405_));
  AOI211_X1 g204(.A(new_n405_), .B(new_n390_), .C1(new_n398_), .C2(new_n402_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n297_), .B(new_n393_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT98), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n397_), .A2(KEYINPUT96), .ZN(new_n409_));
  INV_X1    g208(.A(new_n396_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n402_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n390_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n405_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n403_), .A2(KEYINPUT97), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n394_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT98), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n297_), .A4(new_n393_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G127gat), .B(G134gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G120gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n423_), .ZN(new_n425_));
  AND4_X1   g224(.A1(KEYINPUT94), .A2(new_n258_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(KEYINPUT94), .A2(new_n258_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT4), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n425_), .ZN(new_n429_));
  OR3_X1    g228(.A1(new_n429_), .A2(KEYINPUT4), .A3(new_n258_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n419_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n419_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n426_), .A2(new_n427_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G85gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  OR3_X1    g236(.A1(new_n431_), .A2(new_n433_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT75), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n443_), .B(KEYINPUT30), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(new_n327_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(new_n429_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(G71gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G99gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT31), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n446_), .B(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n408_), .A2(new_n418_), .A3(new_n441_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n385_), .A2(new_n455_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n441_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n439_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n426_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n427_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n461_), .A2(KEYINPUT95), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT95), .B1(new_n461_), .B2(new_n462_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n432_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n437_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n428_), .A2(new_n419_), .A3(new_n430_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT33), .B(new_n437_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n460_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n391_), .A2(new_n470_), .A3(new_n392_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n297_), .B1(new_n458_), .B2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n297_), .A2(new_n440_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(new_n393_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n453_), .B(KEYINPUT78), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n236_), .B1(new_n454_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G57gat), .B(G64gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G71gat), .B(G78gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(KEYINPUT11), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(KEYINPUT11), .ZN(new_n482_));
  INV_X1    g281(.A(new_n480_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n479_), .A2(KEYINPUT11), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n481_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G231gat), .A2(G233gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n214_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n491_));
  XOR2_X1   g290(.A(G127gat), .B(G155gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT16), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G183gat), .B(G211gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(KEYINPUT17), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n490_), .A2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G106gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n450_), .A2(new_n500_), .A3(KEYINPUT66), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT7), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n508_), .A2(new_n450_), .A3(new_n500_), .A4(KEYINPUT66), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n502_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  OR2_X1    g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n511_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT67), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n510_), .A2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT8), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT64), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n524_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n500_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(G92gat), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT9), .ZN(new_n530_));
  AND2_X1   g329(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n512_), .A2(KEYINPUT9), .A3(new_n513_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n507_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n517_), .A2(new_n522_), .B1(new_n528_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n528_), .A2(new_n535_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n538_));
  OAI22_X1  g337(.A1(new_n536_), .A2(new_n224_), .B1(new_n227_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n545_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n539_), .A2(new_n548_), .B1(KEYINPUT36), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n546_), .A2(new_n556_), .A3(new_n547_), .A4(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT37), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n486_), .B(new_n537_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT12), .ZN(new_n562_));
  INV_X1    g361(.A(new_n486_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n538_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(KEYINPUT12), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n565_), .B(new_n566_), .C1(new_n536_), .C2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n564_), .A2(new_n561_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n568_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G120gat), .B(G148gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G176gat), .B(G204gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n570_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(KEYINPUT13), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n577_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n560_), .A2(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n478_), .A2(new_n499_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n440_), .A3(new_n202_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n558_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n454_), .B2(new_n477_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n236_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n580_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n499_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n441_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n584_), .A2(new_n585_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n595_), .A3(new_n596_), .ZN(G1324gat));
  NAND2_X1  g396(.A1(new_n416_), .A2(new_n393_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(G8gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT39), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n583_), .A2(new_n203_), .A3(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT40), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(G1325gat));
  INV_X1    g404(.A(G15gat), .ZN(new_n606_));
  INV_X1    g405(.A(new_n476_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n593_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT99), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT41), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n583_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT100), .Z(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n612_), .A3(new_n614_), .ZN(G1326gat));
  OAI21_X1  g414(.A(G22gat), .B1(new_n594_), .B2(new_n297_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT42), .ZN(new_n617_));
  INV_X1    g416(.A(G22gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n297_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n583_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(G1327gat));
  NOR2_X1   g422(.A1(new_n590_), .A2(new_n499_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n454_), .A2(new_n477_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n626_), .B2(new_n560_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n558_), .B(KEYINPUT37), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT43), .B(new_n628_), .C1(new_n454_), .C2(new_n477_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(KEYINPUT44), .B(new_n624_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(G29gat), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n634_), .A2(new_n635_), .A3(new_n441_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n581_), .A2(new_n499_), .A3(new_n558_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n478_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G29gat), .B1(new_n638_), .B2(new_n440_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n636_), .A2(new_n639_), .ZN(G1328gat));
  INV_X1    g439(.A(G36gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n641_), .A3(new_n598_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT45), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n632_), .A2(new_n598_), .A3(new_n633_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n644_), .A2(new_n645_), .A3(G36gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n644_), .B2(G36gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI221_X1 g449(.A(new_n643_), .B1(KEYINPUT103), .B2(KEYINPUT46), .C1(new_n646_), .C2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  XOR2_X1   g451(.A(KEYINPUT104), .B(G43gat), .Z(new_n653_));
  INV_X1    g452(.A(new_n638_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(new_n476_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n453_), .A2(G43gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n634_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1330gat));
  OAI21_X1  g458(.A(G50gat), .B1(new_n634_), .B2(new_n297_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n297_), .A2(G50gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT106), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(new_n654_), .B2(new_n662_), .ZN(G1331gat));
  AND4_X1   g462(.A1(new_n236_), .A2(new_n588_), .A3(new_n499_), .A4(new_n581_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(G57gat), .A3(new_n440_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT108), .Z(new_n666_));
  AOI21_X1  g465(.A(new_n589_), .B1(new_n454_), .B2(new_n477_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(new_n499_), .A3(new_n581_), .A4(new_n628_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT107), .Z(new_n669_));
  AOI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n440_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n666_), .A2(new_n670_), .ZN(G1332gat));
  INV_X1    g470(.A(G64gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n664_), .B2(new_n598_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT48), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n669_), .A2(new_n672_), .A3(new_n598_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1333gat));
  AOI21_X1  g475(.A(new_n448_), .B1(new_n664_), .B2(new_n607_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT49), .Z(new_n678_));
  NAND3_X1  g477(.A1(new_n669_), .A2(new_n448_), .A3(new_n607_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1334gat));
  INV_X1    g479(.A(G78gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n664_), .B2(new_n619_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT50), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n669_), .A2(new_n681_), .A3(new_n619_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1335gat));
  AND4_X1   g484(.A1(new_n591_), .A2(new_n667_), .A3(new_n581_), .A4(new_n587_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G85gat), .B1(new_n686_), .B2(new_n440_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n627_), .A2(new_n629_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n589_), .A2(new_n499_), .A3(new_n580_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n531_), .A2(new_n532_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n441_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n687_), .B1(new_n691_), .B2(new_n693_), .ZN(G1336gat));
  NAND3_X1  g493(.A1(new_n686_), .A2(new_n529_), .A3(new_n598_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n598_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n697_), .B2(new_n529_), .ZN(G1337gat));
  OAI21_X1  g497(.A(G99gat), .B1(new_n690_), .B2(new_n476_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n686_), .B(new_n453_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g501(.A1(new_n686_), .A2(new_n500_), .A3(new_n619_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n688_), .A2(new_n619_), .A3(new_n689_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT52), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(G106gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n704_), .B2(G106gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g508(.A1(new_n236_), .A2(new_n499_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT109), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n582_), .ZN(new_n712_));
  XOR2_X1   g511(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT54), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n711_), .B(new_n582_), .C1(KEYINPUT110), .C2(new_n715_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT67), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n520_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n537_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n567_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n722_), .A2(new_n723_), .B1(new_n564_), .B2(new_n562_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n724_), .B2(new_n566_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n565_), .B1(new_n536_), .B2(new_n567_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n566_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(KEYINPUT111), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n568_), .A2(KEYINPUT55), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n722_), .A2(new_n723_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n566_), .A4(new_n565_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n729_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n575_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n729_), .B2(new_n734_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n718_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n729_), .A2(new_n734_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT112), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n742_), .A2(KEYINPUT113), .A3(new_n575_), .A4(new_n736_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT56), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n739_), .A2(new_n740_), .A3(new_n743_), .A4(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n570_), .A2(new_n575_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n739_), .A2(new_n744_), .A3(new_n743_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n742_), .A2(KEYINPUT56), .A3(new_n575_), .A4(new_n736_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT114), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n745_), .B(new_n747_), .C1(new_n748_), .C2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n219_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n214_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n220_), .B1(new_n753_), .B2(new_n217_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n232_), .B1(new_n754_), .B2(new_n226_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n235_), .A2(new_n756_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(new_n576_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n751_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n558_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT57), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n746_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n235_), .A2(new_n763_), .A3(new_n756_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n744_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n749_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT58), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n765_), .A2(new_n749_), .ZN(new_n770_));
  OAI211_X1 g569(.A(KEYINPUT115), .B(new_n769_), .C1(new_n770_), .C2(new_n764_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n560_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n587_), .B1(new_n751_), .B2(new_n758_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT57), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n762_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n717_), .B1(new_n591_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n408_), .A2(new_n418_), .A3(new_n453_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n441_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT59), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n761_), .B(new_n587_), .C1(new_n751_), .C2(new_n758_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n772_), .B1(new_n773_), .B2(KEYINPUT57), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n762_), .A2(KEYINPUT117), .A3(new_n772_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n499_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n717_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n778_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n780_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G113gat), .B1(new_n790_), .B2(new_n236_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n776_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n778_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n236_), .A2(G113gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n793_), .B2(new_n794_), .ZN(G1340gat));
  OAI21_X1  g594(.A(G120gat), .B1(new_n790_), .B2(new_n580_), .ZN(new_n796_));
  INV_X1    g595(.A(G120gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n580_), .B2(KEYINPUT60), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(KEYINPUT60), .B2(new_n797_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n796_), .B1(new_n793_), .B2(new_n799_), .ZN(G1341gat));
  NAND2_X1  g599(.A1(new_n499_), .A2(G127gat), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT118), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n780_), .B(new_n802_), .C1(new_n787_), .C2(new_n789_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n792_), .A2(new_n499_), .A3(new_n778_), .ZN(new_n804_));
  INV_X1    g603(.A(G127gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT119), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n803_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1342gat));
  OAI21_X1  g610(.A(G134gat), .B1(new_n790_), .B2(new_n628_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n558_), .A2(G134gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n793_), .B2(new_n813_), .ZN(G1343gat));
  NOR2_X1   g613(.A1(new_n607_), .A2(new_n297_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n416_), .A2(new_n440_), .A3(new_n393_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n775_), .A2(new_n591_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n815_), .B(new_n817_), .C1(new_n818_), .C2(new_n717_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n236_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n580_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n822_), .B(G148gat), .Z(G1345gat));
  XOR2_X1   g622(.A(KEYINPUT61), .B(G155gat), .Z(new_n824_));
  OR3_X1    g623(.A1(new_n819_), .A2(new_n591_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n819_), .B2(new_n591_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1346gat));
  INV_X1    g629(.A(G162gat), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n819_), .A2(new_n831_), .A3(new_n628_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n819_), .B2(new_n558_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n834_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(G1347gat));
  NAND2_X1  g636(.A1(new_n598_), .A2(new_n441_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n476_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n619_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n589_), .B(new_n841_), .C1(new_n786_), .C2(new_n717_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n351_), .B2(new_n347_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT123), .B1(new_n842_), .B2(G169gat), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n844_), .A2(new_n845_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n842_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(G1348gat));
  NOR2_X1   g648(.A1(new_n776_), .A2(new_n619_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(G176gat), .A3(new_n581_), .A4(new_n839_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n581_), .B(new_n841_), .C1(new_n786_), .C2(new_n717_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n852_), .A2(KEYINPUT124), .A3(new_n356_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT124), .B1(new_n852_), .B2(new_n356_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n851_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT125), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n851_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1349gat));
  NAND3_X1  g658(.A1(new_n850_), .A2(new_n499_), .A3(new_n839_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n841_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n787_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n591_), .A2(new_n338_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n860_), .A2(new_n306_), .B1(new_n862_), .B2(new_n863_), .ZN(G1350gat));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n317_), .A3(new_n587_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n787_), .A2(new_n628_), .A3(new_n861_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n307_), .ZN(G1351gat));
  INV_X1    g666(.A(new_n815_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n776_), .A2(new_n868_), .A3(new_n838_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(G197gat), .A3(new_n589_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n871_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G197gat), .B1(new_n869_), .B2(new_n589_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(G1352gat));
  NAND2_X1  g674(.A1(new_n869_), .A2(new_n581_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g676(.A1(new_n792_), .A2(new_n441_), .A3(new_n598_), .A4(new_n815_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n591_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  AND2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n879_), .B2(new_n880_), .ZN(G1354gat));
  AND3_X1   g682(.A1(new_n869_), .A2(G218gat), .A3(new_n560_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n869_), .A2(new_n587_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G218gat), .B1(new_n885_), .B2(KEYINPUT127), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n878_), .B2(new_n558_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n886_), .B2(new_n888_), .ZN(G1355gat));
endmodule


