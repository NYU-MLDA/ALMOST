//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_;
  INV_X1    g000(.A(KEYINPUT8), .ZN(new_n202_));
  XOR2_X1   g001(.A(G85gat), .B(G92gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n205_), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT65), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(KEYINPUT65), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT7), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n202_), .B(new_n203_), .C1(new_n213_), .C2(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT6), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT6), .B1(new_n210_), .B2(new_n211_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT66), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n209_), .A2(new_n221_), .A3(new_n212_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n222_), .A3(new_n215_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n203_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT8), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n223_), .B2(new_n203_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n217_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT12), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(KEYINPUT9), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G106gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT10), .B(G99gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT64), .ZN(new_n235_));
  AOI211_X1 g034(.A(new_n213_), .B(new_n232_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n228_), .A2(new_n229_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n240_));
  XOR2_X1   g039(.A(G71gat), .B(G78gat), .Z(new_n241_));
  OR2_X1    g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n223_), .A2(new_n203_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT67), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT8), .A3(new_n225_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n236_), .B1(new_n249_), .B2(new_n217_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n238_), .B(new_n246_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n228_), .A2(new_n237_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(KEYINPUT69), .A3(KEYINPUT12), .A4(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT70), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n259_), .A3(new_n256_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n256_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n253_), .A2(new_n246_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n250_), .A2(new_n245_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT68), .Z(new_n266_));
  XOR2_X1   g065(.A(G176gat), .B(G204gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G120gat), .B(G148gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT72), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n269_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n261_), .A2(new_n266_), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT13), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n261_), .A2(new_n266_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n272_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT13), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n261_), .A2(new_n266_), .A3(new_n273_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT75), .B(G15gat), .Z(new_n283_));
  INV_X1    g082(.A(G22gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G1gat), .A2(G8gat), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n283_), .A2(new_n284_), .B1(KEYINPUT14), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n284_), .B2(new_n283_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G8gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT76), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n289_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G29gat), .B(G36gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n295_), .B(KEYINPUT15), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n299_), .B2(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G229gat), .A2(G233gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n292_), .B(new_n295_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n304_), .B2(new_n301_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G113gat), .B(G141gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G169gat), .B(G197gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT82), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n305_), .A2(new_n309_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n282_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT102), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT86), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT23), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n319_), .A2(new_n320_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n325_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G169gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT22), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT22), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n320_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT83), .B1(new_n332_), .B2(new_n342_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n326_), .A2(new_n327_), .B1(new_n330_), .B2(new_n329_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n325_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n341_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n320_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G169gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n337_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT83), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n343_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G15gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(G71gat), .B(G99gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT84), .B(G43gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n355_), .A2(new_n361_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n317_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(KEYINPUT86), .A3(new_n362_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G127gat), .B(G134gat), .Z(new_n368_));
  XOR2_X1   g167(.A(G113gat), .B(G120gat), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT85), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G113gat), .B(G120gat), .ZN(new_n373_));
  OR3_X1    g172(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT85), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n373_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n371_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT31), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n365_), .A2(new_n367_), .A3(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n317_), .B(new_n377_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G22gat), .B(G50gat), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n390_));
  OAI22_X1  g189(.A1(new_n390_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G141gat), .A2(G148gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n391_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT87), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(KEYINPUT87), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n389_), .B1(new_n396_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n388_), .B1(new_n386_), .B2(KEYINPUT1), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n388_), .A2(KEYINPUT1), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G141gat), .B(G148gat), .Z(new_n407_));
  AND2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n385_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n390_), .A2(KEYINPUT3), .ZN(new_n410_));
  INV_X1    g209(.A(new_n401_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(new_n399_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n391_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n388_), .B(new_n387_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n406_), .A2(new_n407_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT88), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n409_), .A2(new_n416_), .A3(KEYINPUT29), .ZN(new_n417_));
  XOR2_X1   g216(.A(G211gat), .B(G218gat), .Z(new_n418_));
  INV_X1    g217(.A(KEYINPUT21), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G197gat), .B(G204gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(G211gat), .B(G218gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT21), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n421_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(KEYINPUT21), .A3(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT89), .Z(new_n429_));
  AND2_X1   g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n417_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT90), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n417_), .A2(new_n433_), .A3(new_n430_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT29), .B1(new_n403_), .B2(new_n408_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n428_), .B1(new_n436_), .B2(new_n427_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G78gat), .B(G106gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n384_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n441_), .A3(new_n383_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n409_), .A2(new_n416_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n447_), .A2(KEYINPUT29), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT28), .Z(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n382_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n381_), .A3(new_n450_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n409_), .A2(new_n376_), .A3(new_n416_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n370_), .A2(new_n375_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n414_), .A2(new_n457_), .A3(new_n415_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n414_), .A2(new_n457_), .A3(KEYINPUT94), .A4(new_n415_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n456_), .A2(KEYINPUT4), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT95), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n460_), .A2(new_n461_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT95), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT4), .A4(new_n456_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n409_), .A2(new_n376_), .A3(new_n416_), .A4(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n469_), .B(KEYINPUT97), .Z(new_n470_));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n471_), .B(KEYINPUT96), .Z(new_n472_));
  NAND3_X1  g271(.A1(new_n467_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n464_), .A2(new_n456_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n472_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G1gat), .B(G29gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT0), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n478_), .B(G57gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G85gat), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n473_), .A2(new_n476_), .A3(KEYINPUT101), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n473_), .A2(new_n476_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n483_), .B2(new_n480_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n473_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT101), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n427_), .B1(new_n343_), .B2(new_n352_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT92), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n424_), .A2(new_n426_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n345_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n351_), .B1(new_n345_), .B2(new_n350_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT20), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n344_), .A2(new_n325_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n427_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n491_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT19), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT91), .Z(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT100), .B1(new_n501_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(KEYINPUT20), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n506_), .A2(KEYINPUT92), .B1(new_n499_), .B2(new_n427_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT100), .ZN(new_n508_));
  INV_X1    g307(.A(new_n504_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n497_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n343_), .A2(new_n352_), .A3(new_n427_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n498_), .B(KEYINPUT99), .Z(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT20), .B(new_n512_), .C1(new_n513_), .C2(new_n427_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n503_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G8gat), .B(G36gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT18), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G64gat), .B(G92gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n503_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n512_), .A2(new_n522_), .A3(KEYINPUT20), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n512_), .A2(new_n522_), .A3(KEYINPUT93), .A4(KEYINPUT20), .ZN(new_n526_));
  AOI221_X4 g325(.A(new_n520_), .B1(new_n525_), .B2(new_n526_), .C1(new_n501_), .C2(new_n504_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT27), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n509_), .B1(new_n507_), .B2(new_n497_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n526_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n520_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n501_), .A2(new_n504_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n520_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n521_), .A2(new_n529_), .B1(new_n528_), .B2(new_n537_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n453_), .A2(new_n455_), .B1(new_n488_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n480_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n472_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n474_), .A2(new_n475_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n543_), .A2(new_n536_), .A3(new_n533_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT98), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n473_), .A2(new_n476_), .A3(KEYINPUT33), .A4(new_n480_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT33), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n485_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .A4(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n535_), .B1(new_n534_), .B2(new_n531_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n527_), .A2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n548_), .A2(new_n551_), .A3(new_n546_), .A4(new_n543_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT98), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n535_), .A2(KEYINPUT32), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n530_), .A2(new_n532_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n516_), .B2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n549_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n381_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n453_), .A2(new_n455_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n539_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT35), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT34), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n250_), .A2(new_n296_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT73), .B1(new_n253_), .B2(new_n298_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n568_));
  AOI211_X1 g367(.A(new_n568_), .B(new_n299_), .C1(new_n228_), .C2(new_n237_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n566_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n565_), .A2(new_n562_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT74), .ZN(new_n573_));
  INV_X1    g372(.A(new_n571_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n574_), .B(new_n566_), .C1(new_n567_), .C2(new_n569_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G190gat), .B(G218gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581_));
  INV_X1    g380(.A(new_n579_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n572_), .A2(new_n582_), .A3(new_n575_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n572_), .A2(new_n575_), .ZN(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT36), .B(new_n579_), .C1(new_n585_), .C2(KEYINPUT74), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n561_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT103), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n245_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(new_n292_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT17), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n593_), .B(KEYINPUT69), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n604_));
  NOR2_X1   g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT79), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT79), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(new_n608_), .A3(new_n605_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n602_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT80), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AOI211_X1 g411(.A(KEYINPUT80), .B(new_n602_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n316_), .A2(new_n590_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n488_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n282_), .A2(new_n561_), .A3(new_n313_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n584_), .A2(KEYINPUT37), .A3(new_n586_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT37), .B1(new_n584_), .B2(new_n586_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n607_), .A2(new_n609_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT80), .B1(new_n623_), .B2(new_n602_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT81), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n610_), .A2(new_n611_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT81), .B1(new_n612_), .B2(new_n613_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n622_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n618_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(G1gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n488_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT38), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n617_), .A2(new_n635_), .ZN(G1324gat));
  INV_X1    g435(.A(G8gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n538_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n631_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n615_), .A2(new_n638_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(G8gat), .ZN(new_n642_));
  AOI211_X1 g441(.A(KEYINPUT39), .B(new_n637_), .C1(new_n615_), .C2(new_n638_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(G1325gat));
  OAI21_X1  g445(.A(G15gat), .B1(new_n616_), .B2(new_n381_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT41), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT41), .ZN(new_n649_));
  INV_X1    g448(.A(G15gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n631_), .A2(new_n650_), .A3(new_n382_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(G1326gat));
  NOR2_X1   g451(.A1(new_n451_), .A2(new_n452_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT104), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n284_), .B1(new_n615_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n631_), .A2(new_n284_), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1327gat));
  INV_X1    g458(.A(new_n629_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT37), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n587_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n584_), .A2(new_n586_), .A3(KEYINPUT37), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(KEYINPUT106), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n662_), .A2(new_n666_), .A3(new_n561_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT43), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n622_), .A2(new_n669_), .A3(new_n561_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n660_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n316_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n633_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(KEYINPUT44), .ZN(new_n675_));
  OAI21_X1  g474(.A(G29gat), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n660_), .A2(new_n587_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n618_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n488_), .A2(G29gat), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT107), .Z(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n678_), .B2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n682_), .A2(KEYINPUT108), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(KEYINPUT108), .ZN(new_n684_));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n672_), .A2(KEYINPUT44), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n538_), .B1(new_n672_), .B2(KEYINPUT44), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n618_), .A2(new_n677_), .A3(new_n685_), .A4(new_n638_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT45), .Z(new_n690_));
  OAI211_X1 g489(.A(new_n683_), .B(new_n684_), .C1(new_n688_), .C2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n673_), .A2(new_n638_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G36gat), .B1(new_n692_), .B2(new_n675_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n690_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n693_), .A2(KEYINPUT108), .A3(new_n694_), .A4(new_n682_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n691_), .A2(new_n695_), .ZN(G1329gat));
  NAND3_X1  g495(.A1(new_n673_), .A2(G43gat), .A3(new_n382_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n678_), .A2(new_n381_), .ZN(new_n698_));
  OAI22_X1  g497(.A1(new_n697_), .A2(new_n675_), .B1(G43gat), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g499(.A1(new_n673_), .A2(G50gat), .A3(new_n653_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n618_), .A2(new_n654_), .A3(new_n677_), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n701_), .A2(new_n675_), .B1(G50gat), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT109), .ZN(G1331gat));
  NOR2_X1   g503(.A1(new_n282_), .A2(new_n313_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n561_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(new_n630_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n633_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n282_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n313_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n627_), .A2(new_n628_), .A3(new_n710_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n590_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n633_), .A2(new_n713_), .A3(G57gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n713_), .B2(G57gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n708_), .B1(new_n712_), .B2(new_n715_), .ZN(G1332gat));
  INV_X1    g515(.A(G64gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n707_), .A2(new_n717_), .A3(new_n638_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n712_), .A2(new_n638_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(G64gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT48), .B(new_n717_), .C1(new_n712_), .C2(new_n638_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT111), .ZN(G1333gat));
  INV_X1    g523(.A(G71gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n712_), .B2(new_n382_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT49), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n707_), .A2(new_n725_), .A3(new_n382_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n712_), .B2(new_n654_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT50), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n654_), .A2(new_n730_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT112), .Z(new_n734_));
  NAND2_X1  g533(.A1(new_n707_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1335gat));
  NAND2_X1  g535(.A1(new_n671_), .A2(new_n705_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n488_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n706_), .A2(new_n677_), .ZN(new_n739_));
  INV_X1    g538(.A(G85gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n633_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1336gat));
  OAI21_X1  g541(.A(G92gat), .B1(new_n737_), .B2(new_n538_), .ZN(new_n743_));
  INV_X1    g542(.A(G92gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n744_), .A3(new_n638_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1337gat));
  OAI21_X1  g545(.A(G99gat), .B1(new_n737_), .B2(new_n381_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n739_), .A2(new_n382_), .A3(new_n235_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n233_), .A3(new_n653_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n668_), .A2(new_n670_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n752_), .A2(new_n653_), .A3(new_n629_), .A4(new_n705_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(G106gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G106gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n751_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT114), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n751_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n758_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(new_n614_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n304_), .A2(new_n301_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n308_), .C1(new_n301_), .C2(new_n300_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n310_), .B(new_n768_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n258_), .A2(new_n771_), .A3(new_n260_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n255_), .A2(new_n256_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n771_), .B2(new_n257_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n770_), .B(new_n272_), .C1(new_n772_), .C2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n258_), .A2(new_n771_), .A3(new_n260_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n257_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n773_), .B1(new_n780_), .B2(KEYINPUT55), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n273_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT116), .B1(new_n777_), .B2(KEYINPUT56), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n313_), .B(new_n280_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n769_), .B1(new_n778_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n587_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT57), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n788_), .A3(new_n587_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n280_), .A2(new_n310_), .A3(new_n768_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n791_), .B(KEYINPUT58), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n622_), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n766_), .B1(new_n790_), .B2(new_n798_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n785_), .A2(new_n788_), .A3(new_n587_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n788_), .B1(new_n785_), .B2(new_n587_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n766_), .B(new_n798_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n765_), .B1(new_n799_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n711_), .A2(new_n805_), .A3(new_n282_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n621_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n711_), .B2(new_n282_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT54), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n711_), .A2(new_n282_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT115), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n621_), .A4(new_n806_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n809_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n804_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(G113gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n633_), .A2(new_n538_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n453_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT119), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n816_), .A2(new_n817_), .A3(new_n313_), .A4(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n798_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT118), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n614_), .B1(new_n823_), .B2(new_n802_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n824_), .B2(new_n814_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT59), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n660_), .B1(new_n790_), .B2(new_n798_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n814_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n820_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n826_), .A2(new_n313_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n821_), .B1(new_n831_), .B2(new_n817_), .ZN(G1340gat));
  INV_X1    g631(.A(KEYINPUT60), .ZN(new_n833_));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n709_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n816_), .A2(new_n820_), .A3(new_n836_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n826_), .A2(new_n709_), .A3(new_n830_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n834_), .ZN(G1341gat));
  INV_X1    g638(.A(G127gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n825_), .B2(new_n629_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n765_), .A2(new_n840_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n826_), .A2(new_n830_), .A3(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT120), .B(new_n840_), .C1(new_n825_), .C2(new_n629_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n843_), .A2(new_n845_), .A3(new_n846_), .ZN(G1342gat));
  INV_X1    g646(.A(G134gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n825_), .B2(new_n587_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT121), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n621_), .A2(new_n848_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n826_), .A2(new_n830_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n853_), .B(new_n848_), .C1(new_n825_), .C2(new_n587_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n850_), .A2(new_n852_), .A3(new_n854_), .ZN(G1343gat));
  NOR2_X1   g654(.A1(new_n818_), .A2(new_n455_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT122), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n816_), .A2(new_n313_), .A3(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g658(.A1(new_n816_), .A2(new_n709_), .A3(new_n857_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g660(.A1(new_n816_), .A2(new_n660_), .A3(new_n857_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  AND2_X1   g663(.A1(new_n816_), .A2(new_n857_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n662_), .A2(new_n666_), .A3(G162gat), .ZN(new_n866_));
  INV_X1    g665(.A(new_n587_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n816_), .A2(new_n867_), .A3(new_n857_), .ZN(new_n868_));
  INV_X1    g667(.A(G162gat), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n865_), .A2(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n814_), .A2(new_n827_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n633_), .A2(new_n538_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n381_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n654_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n871_), .A2(new_n710_), .A3(new_n877_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n879_));
  OR3_X1    g678(.A1(new_n878_), .A2(new_n333_), .A3(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n878_), .B2(new_n333_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n348_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n871_), .A2(new_n877_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G176gat), .B1(new_n884_), .B2(new_n709_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n653_), .B1(new_n804_), .B2(new_n815_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n875_), .A2(new_n282_), .A3(new_n337_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n875_), .A2(new_n629_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G183gat), .B1(new_n886_), .B2(new_n890_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n871_), .A2(new_n326_), .A3(new_n765_), .A4(new_n877_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n889_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n326_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n884_), .A2(new_n894_), .A3(new_n614_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n653_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n896_), .B(new_n890_), .C1(new_n824_), .C2(new_n814_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n895_), .B(KEYINPUT124), .C1(G183gat), .C2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n893_), .A2(new_n899_), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n884_), .A2(new_n327_), .A3(new_n867_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n828_), .A2(new_n622_), .A3(new_n876_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n902_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT125), .B1(new_n902_), .B2(G190gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n901_), .B1(new_n903_), .B2(new_n904_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n873_), .A2(new_n455_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n816_), .A2(new_n313_), .A3(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g707(.A1(new_n816_), .A2(new_n906_), .ZN(new_n909_));
  INV_X1    g708(.A(G204gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(KEYINPUT126), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n909_), .A2(new_n709_), .A3(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT126), .B(G204gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n816_), .A2(new_n906_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n282_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n912_), .A2(new_n915_), .ZN(G1353gat));
  XNOR2_X1  g715(.A(KEYINPUT63), .B(G211gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n909_), .A2(new_n614_), .A3(new_n917_), .ZN(new_n918_));
  OAI22_X1  g717(.A1(new_n914_), .A2(new_n765_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1354gat));
  OAI211_X1 g719(.A(new_n867_), .B(new_n906_), .C1(new_n824_), .C2(new_n814_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G218gat), .B1(new_n922_), .B2(KEYINPUT127), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n921_), .A2(new_n924_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n622_), .A2(G218gat), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n923_), .A2(new_n925_), .B1(new_n909_), .B2(new_n926_), .ZN(G1355gat));
endmodule


