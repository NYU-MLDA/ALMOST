//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G127gat), .B(G134gat), .Z(new_n208_));
  XOR2_X1   g007(.A(G113gat), .B(G120gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT81), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n208_), .A2(new_n209_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(KEYINPUT1), .B2(new_n219_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n215_), .A2(new_n224_), .B1(new_n217_), .B2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n227_), .A2(KEYINPUT83), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(KEYINPUT83), .ZN(new_n229_));
  OAI221_X1 g028(.A(new_n226_), .B1(new_n225_), .B2(new_n217_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT84), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n223_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT4), .B1(new_n214_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n213_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n210_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n236_), .B(new_n212_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(new_n233_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n235_), .B1(new_n240_), .B2(KEYINPUT4), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G225gat), .A2(G233gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT89), .Z(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n242_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n240_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n207_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249_));
  INV_X1    g048(.A(new_n247_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n250_), .B(new_n206_), .C1(new_n241_), .C2(new_n244_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n248_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n245_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(KEYINPUT92), .A3(new_n250_), .A4(new_n206_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT27), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT78), .B(G183gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n257_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT23), .ZN(new_n264_));
  INV_X1    g063(.A(G169gat), .ZN(new_n265_));
  INV_X1    g064(.A(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(KEYINPUT24), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(KEYINPUT24), .A3(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n262_), .A2(new_n264_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT79), .B1(new_n265_), .B2(KEYINPUT22), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT22), .B(G169gat), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n266_), .B(new_n273_), .C1(new_n274_), .C2(KEYINPUT79), .ZN(new_n275_));
  INV_X1    g074(.A(G190gat), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n258_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n263_), .B(KEYINPUT23), .Z(new_n278_));
  OAI211_X1 g077(.A(new_n275_), .B(new_n269_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n272_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G197gat), .B(G204gat), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT21), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(KEYINPUT21), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G211gat), .B(G218gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n280_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT20), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT19), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT25), .B(G183gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n257_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n271_), .A2(new_n264_), .A3(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n264_), .B1(G183gat), .B2(G190gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n274_), .A2(new_n266_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n269_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n294_), .B1(new_n301_), .B2(new_n289_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n291_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n280_), .B2(new_n289_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT87), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n289_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT87), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n307_), .B(KEYINPUT20), .C1(new_n280_), .C2(new_n289_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n303_), .B1(new_n309_), .B2(new_n293_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G8gat), .B(G36gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n310_), .A2(new_n316_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n256_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n289_), .B(KEYINPUT86), .C1(new_n233_), .C2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G228gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(G78gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G106gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n322_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n233_), .A2(new_n321_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT28), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n233_), .A2(new_n331_), .A3(new_n321_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT85), .ZN(new_n334_));
  XOR2_X1   g133(.A(G22gat), .B(G50gat), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT85), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n330_), .A2(new_n337_), .A3(new_n332_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n334_), .B2(new_n338_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n328_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n335_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n339_), .A3(new_n327_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n256_), .B1(new_n310_), .B2(new_n316_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n309_), .A2(new_n293_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n291_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT91), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n289_), .B1(new_n301_), .B2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n350_), .B2(new_n301_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n294_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n315_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n347_), .A2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n255_), .A2(new_n320_), .A3(new_n346_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT93), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(KEYINPUT32), .B(new_n316_), .C1(new_n348_), .C2(new_n353_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n310_), .B1(new_n360_), .B2(new_n315_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n252_), .A2(new_n254_), .A3(new_n359_), .A4(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n241_), .A2(new_n246_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n240_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n206_), .B1(new_n365_), .B2(new_n243_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n251_), .A2(new_n363_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n253_), .A2(KEYINPUT33), .A3(new_n250_), .A4(new_n206_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n309_), .A2(new_n293_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n303_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n315_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n367_), .A2(new_n317_), .A3(new_n368_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n362_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n346_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n317_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n377_), .A2(new_n256_), .B1(new_n354_), .B2(new_n347_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n378_), .A2(KEYINPUT93), .A3(new_n255_), .A4(new_n346_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n358_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(G71gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G99gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n280_), .B(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  XNOR2_X1  g186(.A(G15gat), .B(G43gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT80), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n239_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n387_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n320_), .A2(new_n355_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT94), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT94), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n378_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n346_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n255_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(new_n393_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n380_), .A2(new_n393_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G85gat), .B(G92gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n404_), .ZN(new_n406_));
  XOR2_X1   g205(.A(KEYINPUT10), .B(G99gat), .Z(new_n407_));
  INV_X1    g206(.A(G106gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G99gat), .A2(G106gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT6), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n405_), .A2(new_n406_), .A3(new_n409_), .A4(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT8), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT67), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT66), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT66), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT6), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n416_), .A2(new_n418_), .A3(new_n410_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n410_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n414_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n410_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n417_), .A2(KEYINPUT6), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n415_), .A2(KEYINPUT66), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n416_), .A2(new_n418_), .A3(new_n410_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(KEYINPUT67), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT65), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT7), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT7), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT65), .ZN(new_n431_));
  INV_X1    g230(.A(G99gat), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n429_), .A2(new_n431_), .B1(new_n432_), .B2(new_n408_), .ZN(new_n433_));
  AOI211_X1 g232(.A(G99gat), .B(G106gat), .C1(new_n428_), .C2(KEYINPUT7), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n421_), .A2(new_n427_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n402_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n413_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  AOI211_X1 g237(.A(KEYINPUT8), .B(new_n402_), .C1(new_n435_), .C2(new_n411_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n412_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G29gat), .B(G36gat), .Z(new_n441_));
  XOR2_X1   g240(.A(G43gat), .B(G50gat), .Z(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT15), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G232gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT34), .ZN(new_n447_));
  INV_X1    g246(.A(new_n443_), .ZN(new_n448_));
  OAI221_X1 g247(.A(new_n445_), .B1(KEYINPUT35), .B2(new_n447_), .C1(new_n440_), .C2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(KEYINPUT35), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G190gat), .B(G218gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(G134gat), .B(G162gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT71), .B(KEYINPUT72), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT36), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n451_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(new_n457_), .A3(new_n456_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n401_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G230gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(G64gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(G57gat), .ZN(new_n466_));
  INV_X1    g265(.A(G57gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(G64gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(KEYINPUT68), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G57gat), .B(G64gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT68), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT11), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G71gat), .B(G78gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n469_), .A2(KEYINPUT68), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(new_n472_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT11), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT11), .B(new_n475_), .C1(new_n470_), .C2(new_n473_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n440_), .A2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n483_), .B(new_n412_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n464_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(KEYINPUT12), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n440_), .A2(new_n489_), .A3(new_n484_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n486_), .A2(new_n464_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n487_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G120gat), .B(G148gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT5), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G176gat), .B(G204gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n497_), .B(KEYINPUT69), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n493_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n506_));
  OAI22_X1  g305(.A1(new_n499_), .A2(new_n502_), .B1(new_n506_), .B2(KEYINPUT13), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n483_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G231gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G127gat), .B(G155gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT16), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G183gat), .B(G211gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT17), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n523_), .B(KEYINPUT17), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n519_), .A2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT74), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n526_), .B(new_n531_), .C1(new_n519_), .C2(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G169gat), .B(G197gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n516_), .A2(new_n443_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n514_), .B(new_n515_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n448_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n542_), .A3(KEYINPUT76), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT76), .B1(new_n540_), .B2(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n539_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT77), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT77), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n548_), .B(new_n539_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n444_), .A2(new_n541_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(new_n540_), .A3(new_n538_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n537_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n552_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n537_), .ZN(new_n555_));
  AOI211_X1 g354(.A(new_n554_), .B(new_n555_), .C1(new_n547_), .C2(new_n549_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n509_), .A2(new_n534_), .A3(new_n557_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n463_), .A2(KEYINPUT96), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT96), .B1(new_n463_), .B2(new_n558_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(new_n255_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(new_n511_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n401_), .A2(new_n557_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n530_), .A2(new_n532_), .A3(KEYINPUT75), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT75), .B1(new_n530_), .B2(new_n532_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n461_), .B2(KEYINPUT73), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT73), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n459_), .A2(new_n570_), .A3(KEYINPUT37), .A4(new_n460_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n567_), .A2(new_n569_), .A3(new_n508_), .A4(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n564_), .A2(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n574_), .A2(G1gat), .A3(new_n255_), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n563_), .A2(new_n577_), .A3(KEYINPUT97), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT97), .B1(new_n563_), .B2(new_n577_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(G1324gat));
  NAND2_X1  g379(.A1(new_n395_), .A2(new_n397_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n463_), .A2(new_n582_), .A3(new_n558_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(G8gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT98), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT39), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n587_), .A3(G8gat), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n585_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n586_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n582_), .A2(new_n512_), .ZN(new_n591_));
  OAI22_X1  g390(.A1(new_n589_), .A2(new_n590_), .B1(new_n574_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT40), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(G1325gat));
  OR3_X1    g393(.A1(new_n574_), .A2(G15gat), .A3(new_n393_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n392_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n596_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT41), .B1(new_n596_), .B2(G15gat), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n595_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(G1326gat));
  OR3_X1    g400(.A1(new_n574_), .A2(G22gat), .A3(new_n375_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G22gat), .B1(new_n561_), .B2(new_n375_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(KEYINPUT42), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(KEYINPUT42), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n602_), .B1(new_n604_), .B2(new_n605_), .ZN(G1327gat));
  INV_X1    g405(.A(new_n567_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n557_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n508_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n569_), .A2(new_n571_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT43), .B1(new_n401_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n357_), .A2(new_n356_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n392_), .B1(new_n614_), .B2(new_n379_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n581_), .A2(new_n375_), .A3(new_n400_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n613_), .B(new_n610_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n609_), .B1(new_n612_), .B2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(KEYINPUT44), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n380_), .A2(new_n393_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n398_), .A2(new_n400_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n613_), .B1(new_n623_), .B2(new_n610_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n401_), .A2(KEYINPUT43), .A3(new_n611_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT100), .B(new_n620_), .C1(new_n626_), .C2(new_n609_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n618_), .B2(KEYINPUT44), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n619_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(new_n399_), .ZN(new_n631_));
  INV_X1    g430(.A(G29gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n567_), .A2(new_n461_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n564_), .A2(new_n508_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n564_), .A2(KEYINPUT101), .A3(new_n508_), .A4(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n399_), .A2(new_n632_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT102), .ZN(new_n640_));
  OAI22_X1  g439(.A1(new_n631_), .A2(new_n632_), .B1(new_n638_), .B2(new_n640_), .ZN(G1328gat));
  INV_X1    g440(.A(KEYINPUT46), .ZN(new_n642_));
  INV_X1    g441(.A(G36gat), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n636_), .A2(new_n643_), .A3(new_n582_), .A4(new_n637_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT45), .Z(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n630_), .B2(new_n582_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n644_), .B(KEYINPUT45), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n581_), .B(new_n619_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT46), .B(new_n648_), .C1(new_n649_), .C2(new_n643_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(G1329gat));
  NAND3_X1  g450(.A1(new_n630_), .A2(G43gat), .A3(new_n392_), .ZN(new_n652_));
  INV_X1    g451(.A(G43gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(new_n638_), .B2(new_n393_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT47), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT47), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n652_), .A2(new_n657_), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1330gat));
  NOR2_X1   g458(.A1(new_n638_), .A2(new_n375_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(G50gat), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n346_), .A2(G50gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n630_), .B2(new_n662_), .ZN(G1331gat));
  NOR2_X1   g462(.A1(new_n508_), .A2(new_n608_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(new_n567_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n463_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n463_), .A2(KEYINPUT103), .A3(new_n665_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G57gat), .B1(new_n671_), .B2(new_n255_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n401_), .A2(new_n608_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n567_), .A2(new_n569_), .A3(new_n571_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n673_), .A2(new_n509_), .A3(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n467_), .A3(new_n399_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n672_), .A2(new_n676_), .ZN(G1332gat));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n465_), .A3(new_n582_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n668_), .A2(new_n582_), .A3(new_n669_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT48), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G64gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G64gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(G1333gat));
  NAND3_X1  g484(.A1(new_n675_), .A2(new_n382_), .A3(new_n392_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G71gat), .B1(new_n671_), .B2(new_n393_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(KEYINPUT49), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(KEYINPUT49), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(G1334gat));
  NAND2_X1  g489(.A1(new_n346_), .A2(new_n324_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT106), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n675_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G78gat), .B1(new_n671_), .B2(new_n375_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n694_), .A2(new_n696_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n697_), .B2(new_n698_), .ZN(G1335gat));
  NAND3_X1  g498(.A1(new_n673_), .A2(new_n509_), .A3(new_n633_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT107), .ZN(new_n701_));
  INV_X1    g500(.A(G85gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n399_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n607_), .A2(new_n664_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n255_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n703_), .A2(new_n707_), .ZN(G1336gat));
  INV_X1    g507(.A(G92gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n701_), .A2(new_n709_), .A3(new_n582_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G92gat), .B1(new_n706_), .B2(new_n581_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1337gat));
  OR2_X1    g511(.A1(new_n706_), .A2(new_n393_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n392_), .A2(new_n407_), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n713_), .A2(G99gat), .B1(new_n701_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1338gat));
  NAND3_X1  g516(.A1(new_n701_), .A2(new_n408_), .A3(new_n346_), .ZN(new_n718_));
  AOI211_X1 g517(.A(new_n375_), .B(new_n704_), .C1(new_n612_), .C2(new_n617_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT109), .B1(new_n719_), .B2(new_n408_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n722_), .B(G106gat), .C1(new_n706_), .C2(new_n375_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n718_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT53), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n728_), .B(new_n718_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1339gat));
  INV_X1    g529(.A(KEYINPUT59), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT54), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n674_), .A2(new_n732_), .A3(new_n557_), .A4(new_n508_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT54), .B1(new_n572_), .B2(new_n608_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n440_), .A2(new_n489_), .A3(new_n484_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n489_), .B1(new_n440_), .B2(new_n484_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT55), .B(new_n492_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT111), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n491_), .A2(new_n740_), .A3(KEYINPUT55), .A4(new_n492_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n486_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n464_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n492_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n745_));
  XOR2_X1   g544(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n739_), .A2(new_n741_), .A3(new_n744_), .A4(new_n747_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n748_), .A2(KEYINPUT56), .A3(new_n500_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT56), .B1(new_n748_), .B2(new_n500_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(KEYINPUT112), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n500_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(KEYINPUT112), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n498_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n538_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n538_), .B1(new_n516_), .B2(new_n443_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n537_), .B1(new_n551_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n758_), .A2(KEYINPUT113), .A3(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n556_), .A2(new_n765_), .ZN(new_n766_));
  OAI22_X1  g565(.A1(new_n751_), .A2(new_n757_), .B1(new_n503_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT57), .B1(new_n767_), .B2(new_n461_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n503_), .A2(new_n766_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n752_), .A2(new_n753_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n748_), .A2(KEYINPUT56), .A3(new_n500_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n755_), .B1(new_n750_), .B2(KEYINPUT112), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n769_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n462_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n768_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n556_), .A2(new_n765_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n498_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n783_), .B2(KEYINPUT114), .ZN(new_n784_));
  INV_X1    g583(.A(new_n782_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(KEYINPUT114), .C1(new_n750_), .C2(new_n749_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n779_), .B(new_n610_), .C1(new_n784_), .C2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n785_), .B(KEYINPUT58), .C1(new_n750_), .C2(new_n749_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT116), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n749_), .A2(new_n750_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n782_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n780_), .A3(new_n786_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n779_), .B1(new_n795_), .B2(new_n610_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n778_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n735_), .B1(new_n797_), .B2(new_n534_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n398_), .A2(new_n399_), .A3(new_n392_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n731_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n607_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n735_), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n800_), .B(new_n803_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n608_), .A2(G113gat), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n802_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n610_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT115), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n533_), .B1(new_n813_), .B2(new_n778_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT117), .B(new_n801_), .C1(new_n814_), .C2(new_n735_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n608_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(G113gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT118), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n820_), .A3(new_n817_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n808_), .B1(new_n819_), .B2(new_n821_), .ZN(G1340gat));
  NOR3_X1   g621(.A1(new_n802_), .A2(new_n806_), .A3(new_n508_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT120), .B(G120gat), .Z(new_n824_));
  NAND2_X1  g623(.A1(new_n810_), .A2(new_n815_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n508_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(KEYINPUT60), .B2(new_n824_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n823_), .A2(new_n824_), .B1(new_n825_), .B2(new_n827_), .ZN(G1341gat));
  NOR3_X1   g627(.A1(new_n802_), .A2(new_n806_), .A3(new_n534_), .ZN(new_n829_));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n567_), .A2(new_n830_), .ZN(new_n831_));
  OAI22_X1  g630(.A1(new_n829_), .A2(new_n830_), .B1(new_n825_), .B2(new_n831_), .ZN(G1342gat));
  NOR3_X1   g631(.A1(new_n802_), .A2(new_n806_), .A3(new_n611_), .ZN(new_n833_));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n462_), .A2(new_n834_), .ZN(new_n835_));
  OAI22_X1  g634(.A1(new_n833_), .A2(new_n834_), .B1(new_n825_), .B2(new_n835_), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n375_), .A2(new_n392_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n799_), .A2(new_n399_), .A3(new_n581_), .A4(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n557_), .ZN(new_n839_));
  INV_X1    g638(.A(G141gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1344gat));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n508_), .ZN(new_n842_));
  INV_X1    g641(.A(G148gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1345gat));
  NOR2_X1   g643(.A1(new_n838_), .A2(new_n607_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT61), .B(G155gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  OAI21_X1  g646(.A(G162gat), .B1(new_n838_), .B2(new_n611_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n461_), .A2(G162gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n838_), .B2(new_n849_), .ZN(G1347gat));
  NAND2_X1  g649(.A1(new_n582_), .A2(new_n400_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n346_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n567_), .B1(new_n813_), .B2(new_n778_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n608_), .B(new_n852_), .C1(new_n853_), .C2(new_n735_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n804_), .A2(new_n805_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(KEYINPUT121), .A3(new_n608_), .A4(new_n852_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(G169gat), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n857_), .A2(new_n852_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(new_n274_), .A3(new_n608_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n856_), .A2(new_n858_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n863_), .A3(new_n864_), .ZN(G1348gat));
  AOI21_X1  g664(.A(G176gat), .B1(new_n862_), .B2(new_n509_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n798_), .A2(new_n346_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n851_), .A2(new_n266_), .A3(new_n508_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(G1349gat));
  NAND4_X1  g668(.A1(new_n867_), .A2(new_n582_), .A3(new_n400_), .A4(new_n567_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n534_), .A2(new_n295_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n870_), .A2(new_n258_), .B1(new_n862_), .B2(new_n871_), .ZN(G1350gat));
  NAND2_X1  g671(.A1(new_n462_), .A2(new_n257_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n862_), .A2(new_n874_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n862_), .A2(new_n610_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n276_), .ZN(G1351gat));
  NAND2_X1  g676(.A1(new_n837_), .A2(new_n255_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT123), .Z(new_n879_));
  NOR3_X1   g678(.A1(new_n798_), .A2(new_n581_), .A3(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(G197gat), .A3(new_n608_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n883_));
  AOI21_X1  g682(.A(G197gat), .B1(new_n880_), .B2(new_n608_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .ZN(G1352gat));
  AND2_X1   g684(.A1(new_n880_), .A2(new_n509_), .ZN(new_n886_));
  AND2_X1   g685(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n886_), .B2(new_n888_), .ZN(G1353gat));
  NOR3_X1   g689(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n880_), .A2(new_n533_), .A3(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n893_), .B(new_n894_), .Z(G1354gat));
  NAND2_X1  g694(.A1(new_n880_), .A2(new_n462_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT127), .B(G218gat), .Z(new_n897_));
  NOR2_X1   g696(.A1(new_n611_), .A2(new_n897_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n896_), .A2(new_n897_), .B1(new_n880_), .B2(new_n898_), .ZN(G1355gat));
endmodule


