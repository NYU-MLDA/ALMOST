//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT20), .ZN(new_n208_));
  INV_X1    g007(.A(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(KEYINPUT24), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n216_), .A2(KEYINPUT86), .A3(G183gat), .A4(G190gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n217_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n215_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT85), .B1(new_n224_), .B2(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(G183gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT25), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(KEYINPUT84), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(KEYINPUT85), .A3(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G183gat), .ZN(new_n231_));
  INV_X1    g030(.A(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT26), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n229_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n228_), .B(new_n234_), .C1(KEYINPUT84), .C2(new_n227_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n223_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G169gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n210_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT87), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT87), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n240_), .A3(new_n210_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT23), .B1(new_n226_), .B2(new_n232_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(new_n218_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(G169gat), .B2(G176gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n236_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G211gat), .B(G218gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT94), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT94), .ZN(new_n251_));
  INV_X1    g050(.A(G211gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(G218gat), .ZN(new_n253_));
  INV_X1    g052(.A(G218gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(G211gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G197gat), .ZN(new_n258_));
  INV_X1    g057(.A(G204gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT93), .B(G197gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n259_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT95), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n258_), .A2(KEYINPUT93), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n258_), .A2(KEYINPUT93), .ZN(new_n266_));
  OAI21_X1  g065(.A(G204gat), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT95), .A3(new_n260_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n257_), .A2(new_n264_), .A3(KEYINPUT21), .A4(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(new_n259_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT21), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(G197gat), .B2(G204gat), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n250_), .A2(new_n256_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n262_), .A2(new_n271_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n208_), .B1(new_n248_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G226gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT19), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT25), .B(G183gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G190gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n244_), .A2(new_n218_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n282_), .A2(new_n214_), .A3(new_n212_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT98), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n211_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT98), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n283_), .A4(new_n282_), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n213_), .B(KEYINPUT99), .Z(new_n291_));
  OAI211_X1 g090(.A(new_n238_), .B(new_n291_), .C1(new_n222_), .C2(new_n243_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n285_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT95), .B1(new_n267_), .B2(new_n260_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n250_), .A2(new_n256_), .A3(KEYINPUT21), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n296_), .A2(new_n268_), .B1(new_n274_), .B2(new_n273_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n279_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT100), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n285_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n276_), .A2(new_n301_), .A3(KEYINPUT100), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n235_), .A2(new_n223_), .B1(new_n242_), .B2(new_n246_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n208_), .B1(new_n297_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  AOI221_X4 g104(.A(new_n207_), .B1(new_n277_), .B2(new_n298_), .C1(new_n305_), .C2(new_n279_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT27), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT20), .B1(new_n248_), .B2(new_n276_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT100), .B1(new_n276_), .B2(new_n301_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n279_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(new_n302_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n297_), .A2(new_n292_), .A3(new_n284_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n277_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n279_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n206_), .B(KEYINPUT106), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n308_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT107), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n312_), .B1(new_n311_), .B2(new_n302_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n298_), .A2(new_n277_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n207_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n305_), .A2(new_n279_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n206_), .A3(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n321_), .B1(new_n328_), .B2(new_n307_), .ZN(new_n329_));
  AOI211_X1 g128(.A(KEYINPUT107), .B(KEYINPUT27), .C1(new_n325_), .C2(new_n327_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n320_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT90), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT90), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G155gat), .A3(G162gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n337_), .A2(KEYINPUT92), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(KEYINPUT92), .ZN(new_n339_));
  INV_X1    g138(.A(G141gat), .ZN(new_n340_));
  INV_X1    g139(.A(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT3), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(KEYINPUT3), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n343_), .A2(new_n346_), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n338_), .A2(new_n339_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n334_), .A2(new_n336_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT1), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n334_), .A2(new_n336_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n332_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n342_), .A2(new_n344_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n356_), .A2(KEYINPUT91), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT91), .B1(new_n356_), .B2(new_n357_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n350_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n276_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n276_), .A3(new_n363_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n372_), .B(new_n350_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT28), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n356_), .A2(new_n357_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n356_), .A2(KEYINPUT91), .A3(new_n357_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n372_), .A4(new_n350_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n374_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n374_), .B2(new_n381_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n371_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n368_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n374_), .A2(new_n381_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n382_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n374_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n363_), .B1(new_n361_), .B2(new_n276_), .ZN(new_n393_));
  AOI211_X1 g192(.A(new_n364_), .B(new_n297_), .C1(new_n360_), .C2(KEYINPUT29), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n367_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n395_), .A3(new_n371_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n370_), .B1(new_n387_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n369_), .A2(KEYINPUT97), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT97), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n365_), .A2(new_n399_), .A3(new_n366_), .A4(new_n368_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n392_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G127gat), .B(G134gat), .Z(new_n403_));
  XOR2_X1   g202(.A(G113gat), .B(G120gat), .Z(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  NAND2_X1  g204(.A1(new_n360_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n379_), .A2(new_n407_), .A3(new_n350_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n408_), .A3(KEYINPUT4), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n360_), .A2(new_n412_), .A3(new_n405_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n409_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n406_), .A2(new_n408_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT103), .B1(new_n415_), .B2(new_n411_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT103), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n406_), .A2(new_n408_), .A3(new_n417_), .A4(new_n410_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G1gat), .B(G29gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n414_), .A2(new_n416_), .A3(new_n426_), .A4(new_n418_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G71gat), .B(G99gat), .ZN(new_n430_));
  INV_X1    g229(.A(G43gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n303_), .B(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G227gat), .A2(G233gat), .ZN(new_n436_));
  INV_X1    g235(.A(G15gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT30), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n405_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n435_), .B(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n429_), .A2(new_n441_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n331_), .A2(new_n402_), .A3(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n397_), .A2(new_n428_), .A3(new_n401_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n206_), .B1(new_n326_), .B2(new_n323_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n307_), .B1(new_n306_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT107), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n328_), .A2(new_n321_), .A3(new_n307_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n449_), .A3(new_n320_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n416_), .A2(new_n418_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(KEYINPUT104), .A2(KEYINPUT33), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n426_), .A3(new_n414_), .A4(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n306_), .A2(new_n445_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n427_), .A2(new_n452_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n424_), .B1(new_n415_), .B2(new_n410_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT105), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n409_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT105), .B(new_n424_), .C1(new_n415_), .C2(new_n410_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .A4(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n322_), .A2(new_n324_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(new_n464_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n428_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n397_), .A2(new_n401_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n450_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n441_), .B(KEYINPUT89), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n443_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT13), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT72), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n479_), .A2(new_n481_), .A3(KEYINPUT66), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT66), .B1(new_n479_), .B2(new_n481_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT67), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(G99gat), .B2(G106gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT7), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT67), .B1(new_n486_), .B2(KEYINPUT7), .ZN(new_n488_));
  OR2_X1    g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OAI22_X1  g289(.A1(new_n482_), .A2(new_n483_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G85gat), .B(G92gat), .Z(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(KEYINPUT8), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT69), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n479_), .A2(new_n481_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT68), .B1(new_n489_), .B2(new_n484_), .ZN(new_n500_));
  OAI22_X1  g299(.A1(new_n500_), .A2(KEYINPUT7), .B1(new_n489_), .B2(new_n488_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n493_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT8), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n495_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n482_), .A2(new_n483_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT64), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT10), .B(G99gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(G106gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT65), .B(G85gat), .Z(new_n509_));
  INV_X1    g308(.A(G92gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n511_));
  AOI22_X1  g310(.A1(KEYINPUT9), .A2(new_n492_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  OR3_X1    g311(.A1(new_n507_), .A2(new_n506_), .A3(G106gat), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n505_), .A2(new_n508_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n504_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT71), .B(G71gat), .ZN(new_n516_));
  INV_X1    g315(.A(G78gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n515_), .A2(KEYINPUT12), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n480_), .B1(G99gat), .B2(G106gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT69), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n479_), .A2(new_n481_), .A3(new_n496_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n485_), .A2(new_n486_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n534_));
  INV_X1    g333(.A(new_n489_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n484_), .B1(new_n534_), .B2(KEYINPUT68), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n533_), .A2(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n492_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n538_), .A2(KEYINPUT8), .B1(new_n491_), .B2(new_n494_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n514_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n527_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n530_), .B(new_n531_), .C1(new_n487_), .C2(new_n490_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n503_), .B1(new_n542_), .B2(new_n492_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n491_), .A2(new_n494_), .ZN(new_n544_));
  OAI211_X1 g343(.A(KEYINPUT70), .B(new_n514_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n526_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n525_), .B1(new_n546_), .B2(KEYINPUT12), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n541_), .A2(new_n526_), .A3(new_n545_), .ZN(new_n548_));
  INV_X1    g347(.A(G230gat), .ZN(new_n549_));
  INV_X1    g348(.A(G233gat), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n477_), .B1(new_n547_), .B2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n548_), .A2(new_n552_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n545_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT70), .B1(new_n504_), .B2(new_n514_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n524_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT12), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n555_), .A2(new_n560_), .A3(KEYINPUT72), .A4(new_n525_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n548_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n551_), .B1(new_n562_), .B2(new_n546_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G120gat), .B(G148gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n554_), .A2(new_n561_), .A3(new_n563_), .A4(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n569_), .A2(KEYINPUT73), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT73), .B1(new_n569_), .B2(new_n571_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n476_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n571_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT73), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(KEYINPUT73), .A3(new_n571_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(KEYINPUT13), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G29gat), .B(G36gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G43gat), .B(G50gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT15), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G15gat), .B(G22gat), .ZN(new_n585_));
  INV_X1    g384(.A(G1gat), .ZN(new_n586_));
  INV_X1    g385(.A(G8gat), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT14), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G1gat), .B(G8gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n583_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n591_), .B(new_n593_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n595_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT81), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT82), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n596_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(KEYINPUT82), .A3(new_n605_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT83), .Z(new_n612_));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n591_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n526_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT17), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT79), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT80), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n620_), .A2(KEYINPUT17), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n615_), .A2(new_n621_), .A3(new_n625_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n623_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n624_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT34), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT35), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n541_), .A2(new_n583_), .A3(new_n545_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT74), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n541_), .A2(KEYINPUT74), .A3(new_n583_), .A4(new_n545_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n515_), .A2(new_n584_), .B1(new_n633_), .B2(new_n632_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n634_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(new_n636_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n634_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n638_), .A4(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G190gat), .B(G218gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT36), .Z(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT75), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n645_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT77), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n648_), .A2(KEYINPUT36), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n641_), .A2(new_n654_), .A3(new_n644_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT37), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(KEYINPUT76), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT76), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n641_), .A2(new_n654_), .A3(new_n644_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n650_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n662_), .B2(new_n653_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n652_), .A2(new_n659_), .A3(new_n655_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT37), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n629_), .B(new_n658_), .C1(new_n663_), .C2(new_n665_), .ZN(new_n666_));
  NOR4_X1   g465(.A1(new_n475_), .A2(new_n580_), .A3(new_n612_), .A4(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n586_), .A3(new_n428_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT108), .Z(new_n671_));
  OR2_X1    g470(.A1(new_n662_), .A2(KEYINPUT109), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n662_), .A2(KEYINPUT109), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n475_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n611_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n623_), .A2(new_n626_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n580_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n586_), .B1(new_n682_), .B2(new_n428_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n669_), .B2(new_n668_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n671_), .A2(new_n684_), .ZN(G1324gat));
  NAND3_X1  g484(.A1(new_n667_), .A2(new_n587_), .A3(new_n331_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n676_), .A2(new_n680_), .A3(new_n331_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n687_), .A2(new_n688_), .A3(G8gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n687_), .B2(G8gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT111), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n693_), .B(new_n686_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(G1325gat));
  OAI21_X1  g496(.A(G15gat), .B1(new_n681_), .B2(new_n474_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT41), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n667_), .A2(new_n437_), .A3(new_n473_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT112), .ZN(G1326gat));
  INV_X1    g501(.A(G22gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n470_), .B(KEYINPUT113), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n682_), .B2(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT42), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n703_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT114), .Z(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n667_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(G1327gat));
  INV_X1    g509(.A(new_n580_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n662_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n629_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n714_), .A2(new_n475_), .A3(new_n612_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G29gat), .B1(new_n715_), .B2(new_n428_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n658_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n475_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n473_), .B1(new_n450_), .B2(new_n471_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n720_), .B(new_n717_), .C1(new_n721_), .C2(new_n443_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n580_), .A2(new_n677_), .A3(new_n629_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT44), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n428_), .A2(G29gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n716_), .B1(new_n726_), .B2(new_n727_), .ZN(G1328gat));
  INV_X1    g527(.A(G36gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n715_), .A2(new_n729_), .A3(new_n331_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT45), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n726_), .A2(new_n331_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT46), .B(new_n731_), .C1(new_n732_), .C2(new_n729_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n729_), .B1(new_n726_), .B2(new_n331_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n731_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n737_), .ZN(G1329gat));
  AOI21_X1  g537(.A(G43gat), .B1(new_n715_), .B2(new_n473_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n441_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n431_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n726_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g542(.A(G50gat), .B1(new_n715_), .B2(new_n704_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n402_), .A2(G50gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n726_), .B2(new_n745_), .ZN(G1331gat));
  INV_X1    g545(.A(new_n629_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n711_), .A2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n475_), .A2(new_n611_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n718_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(G57gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n428_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n748_), .A2(new_n612_), .A3(new_n676_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(new_n428_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n754_), .B2(new_n751_), .ZN(G1332gat));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n753_), .B2(new_n331_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT48), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n750_), .A2(new_n756_), .A3(new_n331_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n753_), .B2(new_n473_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT49), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n750_), .A2(new_n761_), .A3(new_n473_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1334gat));
  AOI21_X1  g564(.A(new_n517_), .B1(new_n753_), .B2(new_n704_), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n750_), .A2(new_n517_), .A3(new_n704_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1335gat));
  AND2_X1   g569(.A1(new_n580_), .A2(new_n713_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n749_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n428_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n722_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n447_), .A2(new_n448_), .B1(new_n319_), .B2(new_n308_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(new_n429_), .A3(new_n470_), .A4(new_n441_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(new_n444_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n473_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n720_), .B1(new_n779_), .B2(new_n717_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n677_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT116), .B1(new_n580_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n784_), .B(new_n781_), .C1(new_n574_), .C2(new_n579_), .ZN(new_n785_));
  OAI22_X1  g584(.A1(new_n775_), .A2(new_n780_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n428_), .A2(new_n509_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n774_), .B1(new_n787_), .B2(new_n788_), .ZN(G1336gat));
  AOI21_X1  g588(.A(G92gat), .B1(new_n773_), .B2(new_n331_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n331_), .A2(G92gat), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT117), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n787_), .B2(new_n792_), .ZN(G1337gat));
  NOR3_X1   g592(.A1(new_n772_), .A2(new_n740_), .A3(new_n507_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n473_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(G99gat), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT51), .Z(G1338gat));
  OR3_X1    g596(.A1(new_n772_), .A2(G106gat), .A3(new_n470_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n580_), .A2(new_n782_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n784_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n580_), .A2(KEYINPUT116), .A3(new_n782_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n723_), .A2(new_n803_), .A3(KEYINPUT118), .A4(new_n402_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(G106gat), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n786_), .B2(new_n470_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n799_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  AND4_X1   g607(.A1(new_n799_), .A2(new_n807_), .A3(G106gat), .A4(new_n804_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n798_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n798_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  INV_X1    g613(.A(new_n608_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n592_), .A2(new_n594_), .A3(new_n598_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n604_), .B1(new_n597_), .B2(new_n595_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n571_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n554_), .A2(new_n561_), .A3(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n551_), .B1(new_n547_), .B2(new_n562_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n547_), .A2(new_n553_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(KEYINPUT55), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n547_), .A2(new_n553_), .A3(KEYINPUT121), .A4(new_n820_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n821_), .B(new_n822_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n827_), .A2(KEYINPUT56), .A3(new_n568_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n827_), .B2(new_n568_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n819_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT58), .B(new_n819_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n717_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n571_), .A2(KEYINPUT120), .A3(new_n611_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT120), .B1(new_n571_), .B2(new_n611_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n818_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n835_), .B1(new_n841_), .B2(new_n712_), .ZN(new_n842_));
  AOI211_X1 g641(.A(KEYINPUT57), .B(new_n662_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n834_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n747_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n666_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(new_n612_), .A3(new_n579_), .A4(new_n574_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n711_), .A2(new_n612_), .A3(new_n846_), .A4(new_n848_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n845_), .A2(new_n853_), .ZN(new_n854_));
  NOR4_X1   g653(.A1(new_n331_), .A2(new_n402_), .A3(new_n429_), .A4(new_n740_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n844_), .A2(new_n679_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n853_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n860_), .A2(new_n855_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n861_), .B2(new_n856_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n612_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n855_), .ZN(new_n864_));
  OR3_X1    g663(.A1(new_n864_), .A2(G113gat), .A3(new_n677_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1340gat));
  OAI21_X1  g665(.A(G120gat), .B1(new_n862_), .B2(new_n711_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n711_), .A2(KEYINPUT60), .ZN(new_n868_));
  MUX2_X1   g667(.A(new_n868_), .B(KEYINPUT60), .S(G120gat), .Z(new_n869_));
  NAND2_X1  g668(.A1(new_n861_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n870_), .ZN(G1341gat));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n864_), .B2(new_n747_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT122), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n875_), .B(new_n872_), .C1(new_n864_), .C2(new_n747_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n864_), .A2(KEYINPUT59), .B1(new_n854_), .B2(new_n857_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT123), .B(G127gat), .Z(new_n878_));
  NOR2_X1   g677(.A1(new_n679_), .A2(new_n878_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n874_), .A2(new_n876_), .B1(new_n877_), .B2(new_n879_), .ZN(G1342gat));
  OAI21_X1  g679(.A(G134gat), .B1(new_n862_), .B2(new_n718_), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n864_), .A2(G134gat), .A3(new_n674_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1343gat));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n473_), .A2(new_n470_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n859_), .B2(new_n853_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n776_), .A2(new_n428_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n884_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n852_), .B1(new_n679_), .B2(new_n844_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n891_), .A2(KEYINPUT124), .A3(new_n886_), .A4(new_n888_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n611_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G141gat), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n340_), .B(new_n611_), .C1(new_n890_), .C2(new_n892_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1344gat));
  OAI21_X1  g695(.A(new_n580_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G148gat), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n341_), .B(new_n580_), .C1(new_n890_), .C2(new_n892_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1345gat));
  OAI21_X1  g699(.A(new_n629_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n902_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n629_), .B(new_n904_), .C1(new_n890_), .C2(new_n892_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1346gat));
  INV_X1    g705(.A(G162gat), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n907_), .B(new_n675_), .C1(new_n890_), .C2(new_n892_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n887_), .A2(new_n889_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT124), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n887_), .A2(new_n884_), .A3(new_n889_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n718_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n908_), .B1(new_n912_), .B2(new_n907_), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n776_), .A2(new_n428_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n473_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n704_), .A2(new_n915_), .A3(new_n677_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n209_), .B1(new_n854_), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918_));
  OR3_X1    g717(.A1(new_n917_), .A2(new_n918_), .A3(KEYINPUT62), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n854_), .A2(new_n237_), .A3(new_n916_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n917_), .A2(new_n918_), .ZN(new_n921_));
  OAI21_X1  g720(.A(KEYINPUT62), .B1(new_n917_), .B2(new_n918_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n919_), .B(new_n920_), .C1(new_n921_), .C2(new_n922_), .ZN(G1348gat));
  NOR2_X1   g722(.A1(new_n704_), .A2(new_n915_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n854_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G176gat), .B1(new_n925_), .B2(new_n580_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n891_), .A2(new_n402_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n711_), .A2(new_n210_), .A3(new_n915_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1349gat));
  NAND4_X1  g728(.A1(new_n927_), .A2(new_n473_), .A3(new_n629_), .A4(new_n914_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n679_), .A2(new_n280_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n930_), .A2(new_n226_), .B1(new_n925_), .B2(new_n931_), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n854_), .A2(new_n717_), .A3(new_n924_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G190gat), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  AND4_X1   g734(.A1(new_n281_), .A2(new_n854_), .A3(new_n675_), .A4(new_n924_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT126), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n936_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n938_), .A2(new_n939_), .A3(new_n934_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n937_), .A2(new_n940_), .ZN(G1351gat));
  NAND2_X1  g740(.A1(new_n887_), .A2(new_n914_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n677_), .ZN(new_n943_));
  XOR2_X1   g742(.A(KEYINPUT127), .B(G197gat), .Z(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(G1352gat));
  NOR2_X1   g744(.A1(new_n942_), .A2(new_n711_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n259_), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n887_), .A2(new_n678_), .A3(new_n914_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  AND2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n948_), .A2(new_n949_), .A3(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n948_), .B2(new_n949_), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n942_), .B2(new_n718_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n675_), .A2(new_n254_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n942_), .B2(new_n954_), .ZN(G1355gat));
endmodule


