//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_;
  XOR2_X1   g000(.A(KEYINPUT86), .B(KEYINPUT23), .Z(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n202_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT87), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT86), .B(KEYINPUT23), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(new_n205_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n205_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n213_), .B2(new_n208_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n215_), .B1(G169gat), .B2(G176gat), .ZN(new_n216_));
  NOR3_X1   g015(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT85), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(new_n204_), .B2(KEYINPUT26), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n203_), .A2(KEYINPUT25), .ZN(new_n222_));
  OAI221_X1 g021(.A(new_n220_), .B1(new_n221_), .B2(KEYINPUT84), .C1(new_n222_), .C2(KEYINPUT83), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(KEYINPUT83), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(KEYINPUT84), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n203_), .A2(KEYINPUT25), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT85), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .A4(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n214_), .B(new_n218_), .C1(new_n223_), .C2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G169gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n206_), .A2(new_n212_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n210_), .B2(new_n206_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n232_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G43gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G127gat), .B(G134gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G227gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(G15gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT30), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT31), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT2), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G141gat), .ZN(new_n257_));
  INV_X1    g056(.A(G148gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(KEYINPUT89), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n256_), .B1(KEYINPUT3), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(KEYINPUT3), .B2(new_n259_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n261_), .B(new_n262_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n257_), .A2(new_n258_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n264_), .A2(new_n265_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n262_), .B(KEYINPUT1), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n267_), .B(new_n254_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n243_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n243_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(KEYINPUT4), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n277_), .A3(new_n243_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G225gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT97), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G1gat), .B(G29gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n273_), .A2(new_n275_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n282_), .B(new_n288_), .C1(new_n281_), .C2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n281_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n281_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n287_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n253_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G197gat), .B(G204gat), .Z(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT21), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(KEYINPUT21), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n237_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT20), .ZN(new_n308_));
  INV_X1    g107(.A(new_n235_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n214_), .A2(KEYINPUT94), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT94), .B1(new_n214_), .B2(new_n309_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n232_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n234_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n222_), .A2(new_n226_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n221_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(new_n227_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n313_), .B(new_n218_), .C1(new_n314_), .C2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n312_), .A2(new_n305_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n308_), .B1(KEYINPUT95), .B2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n319_), .A2(KEYINPUT95), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT19), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n312_), .A2(new_n318_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(new_n305_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT20), .B1(new_n237_), .B2(new_n306_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n324_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT18), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT96), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n324_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n328_), .A2(new_n325_), .A3(new_n329_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n335_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT27), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n339_), .A2(new_n340_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(KEYINPUT96), .A3(new_n336_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n305_), .A2(KEYINPUT92), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n271_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G233gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(KEYINPUT91), .A2(G228gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(KEYINPUT91), .A2(G228gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n356_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n348_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(KEYINPUT93), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n271_), .A2(KEYINPUT90), .A3(new_n350_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n274_), .B2(KEYINPUT29), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G22gat), .B(G50gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT28), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n361_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n357_), .A2(new_n358_), .A3(new_n348_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OAI22_X1  g171(.A1(new_n360_), .A2(new_n370_), .B1(new_n372_), .B2(new_n359_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n359_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n370_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n374_), .A2(KEYINPUT93), .A3(new_n371_), .A4(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n308_), .B1(new_n327_), .B2(new_n305_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(new_n325_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n330_), .B2(new_n325_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n341_), .B(KEYINPUT27), .C1(new_n380_), .C2(new_n335_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n346_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT100), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n346_), .A2(KEYINPUT100), .A3(new_n377_), .A4(new_n381_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n298_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n335_), .A2(KEYINPUT32), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n296_), .B1(new_n380_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n344_), .B1(KEYINPUT32), .B2(new_n335_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n377_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n295_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n288_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n394_), .B(KEYINPUT99), .C1(new_n281_), .C2(new_n279_), .ZN(new_n395_));
  OAI211_X1 g194(.A(KEYINPUT33), .B(new_n287_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT99), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n279_), .A2(new_n281_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n397_), .B1(new_n398_), .B2(new_n393_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n392_), .A2(new_n395_), .A3(new_n396_), .A4(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n252_), .B1(new_n390_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n377_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n346_), .A2(new_n297_), .A3(new_n381_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n386_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT74), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT12), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G99gat), .A2(G106gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT6), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(G99gat), .A3(G106gat), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n410_), .A2(new_n412_), .A3(KEYINPUT67), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT67), .B1(new_n410_), .B2(new_n412_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT65), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT65), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT10), .ZN(new_n422_));
  INV_X1    g221(.A(G99gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n424_), .B2(new_n417_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n416_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT66), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT9), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT9), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT66), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n428_), .A2(new_n430_), .A3(G85gat), .A4(G92gat), .ZN(new_n431_));
  INV_X1    g230(.A(G85gat), .ZN(new_n432_));
  INV_X1    g231(.A(G92gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G85gat), .A2(G92gat), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n434_), .A2(new_n427_), .A3(KEYINPUT9), .A4(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n431_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n415_), .A2(new_n426_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT68), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT65), .B1(new_n418_), .B2(new_n419_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n424_), .A2(new_n421_), .A3(new_n417_), .ZN(new_n441_));
  AOI21_X1  g240(.A(G106gat), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n431_), .A2(new_n436_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT68), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n415_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n439_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT69), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n410_), .A2(new_n412_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n423_), .A3(new_n416_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n448_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n434_), .A2(new_n435_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT70), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n457_), .A2(KEYINPUT70), .A3(new_n458_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(KEYINPUT8), .A3(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n415_), .A2(new_n454_), .A3(new_n448_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT8), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n458_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n447_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G57gat), .B(G64gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n470_));
  XOR2_X1   g269(.A(G71gat), .B(G78gat), .Z(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n471_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n407_), .B(new_n408_), .C1(new_n468_), .C2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n462_), .A2(KEYINPUT8), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT70), .B1(new_n457_), .B2(new_n458_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n467_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n445_), .B1(new_n444_), .B2(new_n415_), .ZN(new_n480_));
  AND4_X1   g279(.A1(new_n445_), .A2(new_n415_), .A3(new_n426_), .A4(new_n437_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n475_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT74), .B1(new_n483_), .B2(KEYINPUT12), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n476_), .A2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(KEYINPUT73), .B(new_n467_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT73), .B1(new_n463_), .B2(new_n467_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n482_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n475_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT12), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G230gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT64), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n468_), .B2(new_n475_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n485_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n479_), .A2(new_n482_), .A3(new_n475_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT71), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n479_), .A2(new_n482_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n490_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT71), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n479_), .A2(new_n482_), .A3(new_n502_), .A4(new_n475_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT72), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n504_), .A2(new_n505_), .A3(new_n495_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n504_), .B2(new_n495_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n497_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G120gat), .B(G148gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(G176gat), .B(G204gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n508_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n497_), .B(new_n513_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT13), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(KEYINPUT13), .A3(new_n516_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G29gat), .B(G36gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT15), .ZN(new_n527_));
  XOR2_X1   g326(.A(G1gat), .B(G8gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT81), .ZN(new_n529_));
  INV_X1    g328(.A(G22gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n246_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G15gat), .A2(G22gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G1gat), .A2(G8gat), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n531_), .A2(new_n532_), .B1(KEYINPUT14), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n529_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n527_), .A2(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n535_), .A2(new_n526_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n535_), .B(new_n526_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n540_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n521_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n406_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT36), .Z(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT34), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT35), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n479_), .A2(new_n482_), .A3(new_n526_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT78), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT78), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n479_), .A2(new_n482_), .A3(new_n564_), .A4(new_n526_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n561_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n489_), .A2(new_n527_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n560_), .A2(KEYINPUT35), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n558_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n568_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n571_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n558_), .B(KEYINPUT79), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n578_), .B1(new_n582_), .B2(new_n577_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT80), .B1(new_n579_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT80), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n571_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n582_), .A2(new_n577_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n585_), .B(new_n586_), .C1(new_n587_), .C2(new_n578_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n475_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n535_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G127gat), .B(G155gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n596_), .A2(new_n597_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n592_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT82), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT82), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n599_), .A2(new_n604_), .A3(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n589_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n554_), .A2(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n609_), .A2(G1gat), .A3(new_n297_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT38), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n571_), .A2(new_n577_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n406_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n553_), .A2(new_n607_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n297_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n610_), .A2(KEYINPUT38), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n617_), .A3(new_n618_), .ZN(G1324gat));
  NAND2_X1  g418(.A1(new_n346_), .A2(new_n381_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n609_), .A2(G8gat), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G8gat), .B1(new_n616_), .B2(new_n621_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(G8gat), .B(new_n624_), .C1(new_n616_), .C2(new_n621_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n622_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n628_), .B(new_n629_), .Z(G1325gat));
  OAI21_X1  g429(.A(G15gat), .B1(new_n616_), .B2(new_n252_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT41), .Z(new_n632_));
  INV_X1    g431(.A(new_n609_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n246_), .A3(new_n253_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n616_), .B2(new_n377_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT42), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n530_), .A3(new_n403_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n553_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n612_), .A2(new_n606_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n640_), .B(new_n641_), .C1(new_n386_), .C2(new_n405_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n296_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n589_), .B1(new_n386_), .B2(new_n405_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT43), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n647_), .B(new_n589_), .C1(new_n386_), .C2(new_n405_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n553_), .A2(new_n606_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n650_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n296_), .A2(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n644_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n653_), .A2(new_n620_), .A3(new_n654_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G36gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n621_), .A2(G36gat), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n642_), .A2(KEYINPUT45), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT45), .B1(new_n642_), .B2(new_n665_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n658_), .A2(new_n659_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n661_), .B1(new_n663_), .B2(new_n671_), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n660_), .B(new_n670_), .C1(new_n662_), .C2(G36gat), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1329gat));
  NAND4_X1  g473(.A1(new_n653_), .A2(G43gat), .A3(new_n253_), .A4(new_n654_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n642_), .A2(new_n252_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(G43gat), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n675_), .B(new_n678_), .C1(G43gat), .C2(new_n676_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1330gat));
  AOI21_X1  g481(.A(G50gat), .B1(new_n643_), .B2(new_n403_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n403_), .A2(G50gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n655_), .B2(new_n684_), .ZN(G1331gat));
  INV_X1    g484(.A(new_n521_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n614_), .A2(new_n606_), .A3(new_n551_), .A4(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G57gat), .B1(new_n687_), .B2(new_n297_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n406_), .A2(new_n552_), .A3(new_n521_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n608_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n297_), .A2(G57gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT105), .ZN(G1332gat));
  OAI21_X1  g492(.A(G64gat), .B1(new_n687_), .B2(new_n621_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT48), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n621_), .A2(G64gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n690_), .B2(new_n696_), .ZN(G1333gat));
  OAI21_X1  g496(.A(G71gat), .B1(new_n687_), .B2(new_n252_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT49), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n252_), .A2(G71gat), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT106), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n690_), .B2(new_n701_), .ZN(G1334gat));
  OAI21_X1  g501(.A(G78gat), .B1(new_n687_), .B2(new_n377_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n377_), .A2(G78gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n690_), .B2(new_n706_), .ZN(G1335gat));
  NAND2_X1  g506(.A1(new_n689_), .A2(new_n641_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n432_), .A3(new_n296_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n686_), .A2(new_n607_), .A3(new_n551_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT108), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n713_), .A2(new_n714_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n297_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n710_), .B1(new_n717_), .B2(new_n432_), .ZN(G1336gat));
  NAND3_X1  g517(.A1(new_n709_), .A2(new_n433_), .A3(new_n620_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n715_), .A2(new_n716_), .A3(new_n621_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n433_), .ZN(G1337gat));
  OAI211_X1 g520(.A(new_n709_), .B(new_n253_), .C1(new_n420_), .C2(new_n425_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n713_), .A2(new_n253_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(G99gat), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT110), .B(new_n423_), .C1(new_n713_), .C2(new_n253_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT51), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(new_n722_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1338gat));
  NAND3_X1  g530(.A1(new_n709_), .A2(new_n416_), .A3(new_n403_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n713_), .A2(new_n403_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G106gat), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT52), .B(new_n416_), .C1(new_n713_), .C2(new_n403_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n732_), .B(new_n738_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1339gat));
  AOI211_X1 g541(.A(new_n297_), .B(new_n252_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT59), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n606_), .A2(new_n551_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n519_), .A2(new_n520_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT112), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n584_), .A2(new_n588_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n519_), .A2(new_n750_), .A3(new_n520_), .A4(new_n746_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n748_), .A2(new_n749_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT113), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n747_), .A2(KEYINPUT112), .B1(new_n584_), .B2(new_n588_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n759_), .A3(new_n751_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n755_), .A2(new_n756_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n756_), .B1(new_n755_), .B2(new_n760_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n543_), .A2(new_n539_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n547_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT116), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n538_), .A2(new_n539_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n537_), .B2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(KEYINPUT116), .A3(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n517_), .A2(new_n548_), .A3(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n552_), .A2(new_n516_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n499_), .A2(new_n503_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n485_), .A2(new_n493_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n495_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n497_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n485_), .A2(KEYINPUT55), .A3(new_n493_), .A4(new_n496_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT115), .B1(new_n779_), .B2(new_n514_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n772_), .B1(new_n780_), .B2(KEYINPUT56), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  AOI211_X1 g581(.A(KEYINPUT115), .B(new_n782_), .C1(new_n779_), .C2(new_n514_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n771_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT57), .A3(new_n612_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(KEYINPUT118), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n779_), .A2(new_n514_), .A3(new_n787_), .A4(new_n788_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n770_), .A2(new_n548_), .A3(new_n516_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n776_), .A2(new_n497_), .B1(new_n774_), .B2(new_n495_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n513_), .B1(new_n791_), .B2(new_n778_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n789_), .B(new_n790_), .C1(new_n792_), .C2(new_n787_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n779_), .A2(new_n514_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n786_), .A3(KEYINPUT56), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n797_), .A2(KEYINPUT58), .A3(new_n789_), .A4(new_n790_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n589_), .A2(new_n795_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n785_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT57), .B1(new_n784_), .B2(new_n612_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n607_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n745_), .B1(new_n763_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n784_), .A2(new_n612_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT117), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(new_n800_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n801_), .A2(KEYINPUT117), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n606_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n760_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n757_), .A2(new_n751_), .B1(KEYINPUT113), .B2(new_n753_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT114), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n755_), .A2(new_n756_), .A3(new_n760_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT119), .B1(new_n809_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n808_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n785_), .B(new_n799_), .C1(new_n801_), .C2(KEYINPUT117), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n607_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n763_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(new_n820_), .A3(new_n743_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n803_), .B1(new_n821_), .B2(KEYINPUT59), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n822_), .A2(new_n552_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n552_), .A2(new_n824_), .ZN(new_n825_));
  OAI22_X1  g624(.A1(new_n823_), .A2(new_n824_), .B1(new_n821_), .B2(new_n825_), .ZN(G1340gat));
  AND2_X1   g625(.A1(new_n822_), .A2(new_n686_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT120), .B(G120gat), .Z(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n521_), .B2(KEYINPUT60), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(KEYINPUT60), .B2(new_n828_), .ZN(new_n830_));
  OAI22_X1  g629(.A1(new_n827_), .A2(new_n828_), .B1(new_n821_), .B2(new_n830_), .ZN(G1341gat));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833_));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n607_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n803_), .B(new_n836_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n815_), .A2(new_n820_), .A3(new_n743_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G127gat), .B1(new_n838_), .B2(new_n606_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n832_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n803_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n836_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(new_n842_), .C1(new_n838_), .C2(new_n744_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n834_), .B1(new_n821_), .B2(new_n607_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(KEYINPUT122), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n845_), .ZN(G1342gat));
  INV_X1    g645(.A(G134gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n821_), .B2(new_n612_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT123), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n850_), .B(new_n847_), .C1(new_n821_), .C2(new_n612_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n749_), .A2(new_n847_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n849_), .A2(new_n851_), .B1(new_n822_), .B2(new_n852_), .ZN(G1343gat));
  AND2_X1   g652(.A1(new_n815_), .A2(new_n820_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n403_), .A2(new_n252_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n620_), .A2(new_n855_), .A3(new_n297_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n552_), .A3(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g657(.A1(new_n854_), .A2(new_n686_), .A3(new_n856_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g659(.A1(new_n854_), .A2(new_n606_), .A3(new_n856_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  NAND2_X1  g662(.A1(new_n854_), .A2(new_n856_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G162gat), .B1(new_n864_), .B2(new_n749_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n612_), .A2(G162gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n864_), .B2(new_n866_), .ZN(G1347gat));
  AOI21_X1  g666(.A(new_n403_), .B1(new_n763_), .B2(new_n802_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n621_), .A2(new_n298_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n552_), .A3(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n871_));
  AND4_X1   g670(.A1(KEYINPUT125), .A2(new_n870_), .A3(G169gat), .A4(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(G169gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n871_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n870_), .A2(new_n876_), .B1(KEYINPUT125), .B2(new_n871_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT22), .B(G169gat), .Z(new_n878_));
  OAI22_X1  g677(.A1(new_n872_), .A2(new_n877_), .B1(new_n870_), .B2(new_n878_), .ZN(G1348gat));
  NAND2_X1  g678(.A1(new_n868_), .A2(new_n869_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n521_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(G176gat), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n854_), .A2(new_n377_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n869_), .A2(G176gat), .A3(new_n686_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n882_), .B1(new_n883_), .B2(new_n885_), .ZN(G1349gat));
  NOR3_X1   g685(.A1(new_n621_), .A2(new_n607_), .A3(new_n298_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n868_), .A2(new_n314_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n883_), .A2(new_n887_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n203_), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n868_), .A2(new_n589_), .A3(new_n869_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G190gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n613_), .A2(new_n316_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n880_), .B2(new_n893_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT126), .ZN(G1351gat));
  NOR3_X1   g694(.A1(new_n621_), .A2(new_n296_), .A3(new_n855_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n854_), .A2(new_n552_), .A3(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g697(.A1(new_n854_), .A2(new_n686_), .A3(new_n896_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g699(.A(new_n607_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n854_), .A2(new_n896_), .A3(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n902_), .B(new_n903_), .Z(G1354gat));
  AND2_X1   g703(.A1(new_n854_), .A2(new_n896_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n613_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT127), .B(G218gat), .Z(new_n907_));
  NOR2_X1   g706(.A1(new_n749_), .A2(new_n907_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n906_), .A2(new_n907_), .B1(new_n905_), .B2(new_n908_), .ZN(G1355gat));
endmodule


