//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n203_), .A2(new_n204_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT8), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n211_), .A2(new_n212_), .B1(new_n213_), .B2(KEYINPUT66), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(KEYINPUT66), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT7), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n214_), .B1(new_n215_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G85gat), .ZN(new_n227_));
  INV_X1    g026(.A(G92gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n210_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n210_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n222_), .A2(new_n224_), .A3(KEYINPUT65), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT65), .B1(new_n222_), .B2(new_n224_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n220_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n233_), .B1(new_n236_), .B2(KEYINPUT67), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n220_), .B(new_n238_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n232_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n234_), .A2(new_n235_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT9), .ZN(new_n242_));
  INV_X1    g041(.A(new_n230_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n242_), .B(new_n229_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n229_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n230_), .ZN(new_n246_));
  OR2_X1    g045(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n212_), .A3(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n209_), .B1(new_n240_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n219_), .A2(new_n215_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n214_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT67), .B1(new_n241_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n233_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n239_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n232_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n234_), .A2(new_n235_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n246_), .A2(new_n249_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n262_), .A2(KEYINPUT68), .A3(new_n245_), .A4(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(new_n241_), .B2(new_n250_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n261_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n209_), .A2(KEYINPUT12), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n252_), .A2(new_n253_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G230gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n251_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n209_), .ZN(new_n275_));
  AOI211_X1 g074(.A(KEYINPUT69), .B(new_n273_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n277_));
  INV_X1    g076(.A(new_n251_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n261_), .A2(new_n278_), .A3(new_n275_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n279_), .B2(new_n272_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n271_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n240_), .A2(new_n251_), .A3(new_n209_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n275_), .B1(new_n261_), .B2(new_n278_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n273_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT5), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G176gat), .B(G204gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(new_n284_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT70), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n281_), .A2(new_n292_), .A3(new_n284_), .A4(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n281_), .A2(new_n284_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n288_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT13), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(KEYINPUT13), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n297_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G231gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n209_), .B(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G1gat), .B(G8gat), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G15gat), .B(G22gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311_));
  INV_X1    g110(.A(G1gat), .ZN(new_n312_));
  INV_X1    g111(.A(G8gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT14), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n311_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n309_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n308_), .A3(new_n315_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n307_), .B(new_n321_), .Z(new_n322_));
  XNOR2_X1  g121(.A(G127gat), .B(G155gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT16), .ZN(new_n324_));
  XOR2_X1   g123(.A(G183gat), .B(G211gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT17), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n326_), .A2(new_n327_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n322_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n328_), .B2(new_n322_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT78), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G229gat), .A2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G43gat), .B(G50gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G36gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G29gat), .ZN(new_n339_));
  INV_X1    g138(.A(G29gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G36gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT73), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT73), .B1(new_n339_), .B2(new_n341_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n337_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n341_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(new_n342_), .A3(new_n336_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n350_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n335_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n321_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(KEYINPUT80), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n334_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT15), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n350_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n345_), .A2(new_n349_), .A3(KEYINPUT15), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n321_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n334_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G113gat), .B(G141gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G169gat), .B(G197gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  NOR2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n368_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n358_), .A2(new_n364_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n353_), .A2(new_n357_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n334_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n364_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n368_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(KEYINPUT81), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n369_), .B1(new_n373_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n373_), .A2(new_n380_), .A3(new_n369_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n305_), .A2(new_n333_), .A3(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G190gat), .B(G218gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G134gat), .B(G162gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT36), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n360_), .A2(new_n361_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT75), .B1(new_n268_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT74), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n274_), .A2(new_n350_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G232gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .A4(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n397_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT35), .B1(new_n392_), .B2(new_n394_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n390_), .B(new_n399_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n392_), .A2(new_n394_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n400_), .B(new_n397_), .C1(new_n406_), .C2(KEYINPUT35), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n407_), .A2(KEYINPUT76), .A3(new_n390_), .A4(new_n399_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n399_), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n389_), .B(KEYINPUT36), .Z(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT88), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT25), .B(G183gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT26), .B(G190gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(G169gat), .B2(G176gat), .ZN(new_n422_));
  NOR3_X1   g221(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT23), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n416_), .A2(new_n417_), .A3(KEYINPUT83), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n420_), .A2(new_n424_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(G183gat), .B2(G190gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G169gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT86), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n428_), .A2(KEYINPUT30), .A3(new_n432_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT31), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n436_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G127gat), .B(G134gat), .Z(new_n442_));
  XOR2_X1   g241(.A(G113gat), .B(G120gat), .Z(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G127gat), .B(G134gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G113gat), .B(G120gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT87), .B1(new_n444_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(KEYINPUT87), .A3(new_n447_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(G15gat), .ZN(new_n452_));
  INV_X1    g251(.A(G43gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G15gat), .A2(G43gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G71gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(KEYINPUT84), .A3(new_n455_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n463_));
  OAI21_X1  g262(.A(G99gat), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n458_), .A2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(G71gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n211_), .A3(new_n461_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n468_), .B(KEYINPUT85), .Z(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n464_), .A2(new_n467_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n441_), .A2(new_n451_), .A3(new_n470_), .A4(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n451_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n470_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n475_), .B1(new_n476_), .B2(new_n440_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n438_), .A2(KEYINPUT31), .ZN(new_n478_));
  AND4_X1   g277(.A1(new_n439_), .A2(new_n474_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n474_), .A2(new_n477_), .B1(new_n478_), .B2(new_n439_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n415_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n477_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n439_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n474_), .A2(new_n477_), .A3(new_n439_), .A4(new_n478_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(KEYINPUT88), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G211gat), .B(G218gat), .Z(new_n488_));
  OR2_X1    g287(.A1(G197gat), .A2(G204gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT91), .B(G197gat), .ZN(new_n490_));
  INV_X1    g289(.A(G204gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT21), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n488_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(G197gat), .B2(G204gat), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n495_), .A2(KEYINPUT92), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT92), .B1(new_n495_), .B2(new_n496_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n488_), .A2(KEYINPUT21), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(new_n492_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT93), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n504_), .A3(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G228gat), .A2(G233gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT90), .Z(new_n507_));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n508_));
  INV_X1    g307(.A(G141gat), .ZN(new_n509_));
  INV_X1    g308(.A(G148gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G141gat), .A2(G148gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT2), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n511_), .A2(new_n514_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G155gat), .ZN(new_n518_));
  INV_X1    g317(.A(G162gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT89), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(G155gat), .B2(G162gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G155gat), .A2(G162gat), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n517_), .A2(new_n520_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT1), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT1), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(G155gat), .A3(G162gat), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n525_), .A2(new_n520_), .A3(new_n522_), .A4(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n509_), .A2(new_n510_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n512_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT29), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n503_), .A2(new_n505_), .A3(new_n507_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n502_), .A2(new_n532_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n507_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G78gat), .B(G106gat), .Z(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n533_), .A2(new_n540_), .A3(new_n536_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n531_), .A2(KEYINPUT29), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT28), .ZN(new_n544_));
  XOR2_X1   g343(.A(G22gat), .B(G50gat), .Z(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n539_), .A2(new_n546_), .A3(new_n547_), .A4(new_n541_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n487_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n503_), .A2(new_n505_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(new_n432_), .A3(new_n428_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G226gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT19), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n432_), .B(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n424_), .A2(new_n418_), .A3(new_n426_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n558_), .B1(new_n562_), .B2(new_n502_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n557_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n432_), .A2(new_n561_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT20), .B1(new_n502_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n503_), .A2(new_n433_), .A3(new_n505_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT95), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n503_), .A2(new_n569_), .A3(new_n433_), .A4(new_n505_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n566_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n564_), .B1(new_n571_), .B2(new_n557_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G8gat), .B(G36gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(G64gat), .B(G92gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT32), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n572_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT101), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n572_), .A2(new_n583_), .A3(new_n580_), .ZN(new_n584_));
  OAI211_X1 g383(.A(KEYINPUT20), .B(new_n557_), .C1(new_n562_), .C2(new_n502_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n557_), .B1(new_n554_), .B2(new_n563_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n579_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G1gat), .B(G29gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G85gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT0), .B(G57gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G225gat), .A2(G233gat), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n444_), .A2(KEYINPUT87), .A3(new_n447_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n531_), .B1(new_n597_), .B2(new_n448_), .ZN(new_n598_));
  OR2_X1    g397(.A1(KEYINPUT99), .A2(KEYINPUT4), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(KEYINPUT98), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n444_), .A2(new_n447_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n531_), .B(new_n605_), .C1(new_n597_), .C2(new_n448_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n451_), .A2(KEYINPUT99), .A3(new_n531_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n596_), .B(new_n601_), .C1(new_n609_), .C2(KEYINPUT4), .ZN(new_n610_));
  INV_X1    g409(.A(new_n596_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n595_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n608_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n606_), .A2(new_n604_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n615_), .B2(new_n602_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT4), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n611_), .B(new_n600_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n612_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n594_), .A3(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n613_), .A2(KEYINPUT102), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n622_), .B(new_n595_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n590_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n607_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n594_), .B1(new_n626_), .B2(new_n611_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n601_), .B1(new_n609_), .B2(KEYINPUT4), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n596_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n628_), .B2(new_n596_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n618_), .A2(KEYINPUT33), .A3(new_n594_), .A4(new_n619_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n620_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n588_), .A2(KEYINPUT97), .A3(new_n578_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n568_), .A2(new_n570_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n585_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n554_), .A2(new_n563_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n556_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n642_), .A3(new_n578_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n577_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n636_), .B1(new_n637_), .B2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n552_), .B1(new_n625_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n624_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n621_), .A2(KEYINPUT103), .A3(new_n623_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT27), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n646_), .A2(new_n653_), .A3(new_n637_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n572_), .A2(new_n577_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(KEYINPUT27), .A3(new_n643_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n481_), .A2(new_n551_), .A3(new_n486_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n549_), .B(new_n550_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n652_), .A2(new_n657_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n414_), .B1(new_n648_), .B2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n386_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n652_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n304_), .B(KEYINPUT72), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT37), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n413_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n409_), .A2(KEYINPUT37), .A3(new_n412_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n333_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n668_), .A2(KEYINPUT79), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT79), .ZN(new_n675_));
  INV_X1    g474(.A(new_n673_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n667_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n648_), .A2(new_n661_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n674_), .A2(new_n677_), .A3(new_n384_), .A4(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n652_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n312_), .A3(new_n680_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT104), .A3(new_n666_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT104), .B1(new_n681_), .B2(new_n666_), .ZN(new_n683_));
  OAI221_X1 g482(.A(new_n665_), .B1(new_n666_), .B2(new_n681_), .C1(new_n682_), .C2(new_n683_), .ZN(G1324gat));
  OAI21_X1  g483(.A(G8gat), .B1(new_n664_), .B2(new_n657_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT39), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n654_), .A2(new_n656_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n679_), .A2(new_n313_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n689_), .B(new_n691_), .ZN(G1325gat));
  AOI21_X1  g491(.A(new_n452_), .B1(new_n663_), .B2(new_n487_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT41), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n679_), .A2(new_n452_), .A3(new_n487_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1326gat));
  INV_X1    g495(.A(G22gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n663_), .B2(new_n551_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT106), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(KEYINPUT42), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(KEYINPUT42), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n679_), .A2(new_n697_), .A3(new_n551_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(G1327gat));
  NAND3_X1  g502(.A1(new_n304_), .A2(new_n333_), .A3(new_n384_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  AOI211_X1 g507(.A(new_n707_), .B(new_n708_), .C1(new_n678_), .C2(new_n672_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n621_), .A2(KEYINPUT103), .A3(new_n623_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT103), .B1(new_n621_), .B2(new_n623_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n660_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(new_n687_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n487_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n551_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n646_), .A2(new_n637_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n717_), .A2(new_n632_), .A3(new_n633_), .A4(new_n635_), .ZN(new_n718_));
  AOI22_X1  g517(.A1(new_n581_), .A2(KEYINPUT101), .B1(new_n588_), .B2(new_n579_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n719_), .A2(new_n623_), .A3(new_n621_), .A4(new_n584_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n716_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n672_), .B1(new_n713_), .B2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT43), .B1(new_n722_), .B2(KEYINPUT108), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n706_), .B1(new_n709_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n706_), .B(KEYINPUT44), .C1(new_n709_), .C2(new_n723_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(G29gat), .A3(new_n680_), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n413_), .B(new_n332_), .C1(new_n648_), .C2(new_n661_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n305_), .A2(new_n385_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n340_), .B1(new_n732_), .B2(new_n652_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(G1328gat));
  INV_X1    g535(.A(new_n732_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n687_), .A2(KEYINPUT111), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n687_), .A2(KEYINPUT111), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n737_), .A2(new_n338_), .A3(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT45), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n726_), .A2(new_n687_), .A3(new_n727_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(G36gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G36gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT46), .B(new_n743_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1329gat));
  NOR2_X1   g551(.A1(new_n479_), .A2(new_n480_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n728_), .A2(G43gat), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n453_), .B1(new_n732_), .B2(new_n714_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g557(.A(G50gat), .B1(new_n737_), .B2(new_n551_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n551_), .A2(G50gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n728_), .B2(new_n760_), .ZN(G1331gat));
  AND4_X1   g560(.A1(new_n673_), .A2(new_n678_), .A3(new_n305_), .A4(new_n385_), .ZN(new_n762_));
  INV_X1    g561(.A(G57gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n680_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n668_), .A2(new_n384_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(new_n332_), .A3(new_n662_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(new_n680_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n764_), .B1(new_n767_), .B2(new_n763_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT112), .Z(G1332gat));
  INV_X1    g568(.A(G64gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n766_), .B2(new_n741_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT48), .Z(new_n772_));
  NAND3_X1  g571(.A1(new_n762_), .A2(new_n770_), .A3(new_n741_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1333gat));
  AOI21_X1  g573(.A(new_n459_), .B1(new_n766_), .B2(new_n487_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT49), .Z(new_n776_));
  NAND3_X1  g575(.A1(new_n762_), .A2(new_n459_), .A3(new_n487_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1334gat));
  INV_X1    g577(.A(G78gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n766_), .B2(new_n551_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT50), .Z(new_n781_));
  NAND3_X1  g580(.A1(new_n762_), .A2(new_n779_), .A3(new_n551_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1335gat));
  OR2_X1    g582(.A1(new_n709_), .A2(new_n723_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n304_), .A2(new_n332_), .A3(new_n384_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G85gat), .B1(new_n786_), .B2(new_n652_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n765_), .A2(new_n730_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(new_n227_), .A3(new_n680_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1336gat));
  OAI21_X1  g589(.A(G92gat), .B1(new_n786_), .B2(new_n740_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(new_n228_), .A3(new_n687_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1337gat));
  NAND4_X1  g592(.A1(new_n788_), .A2(new_n247_), .A3(new_n248_), .A4(new_n754_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n784_), .A2(new_n487_), .A3(new_n785_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n795_), .A2(KEYINPUT113), .A3(G99gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT113), .B1(new_n795_), .B2(G99gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n788_), .A2(new_n212_), .A3(new_n551_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n784_), .A2(new_n551_), .A3(new_n785_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G106gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT53), .ZN(G1339gat));
  OR3_X1    g605(.A1(new_n652_), .A2(new_n687_), .A3(new_n659_), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT117), .Z(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR4_X1   g608(.A1(new_n305_), .A2(new_n672_), .A3(new_n333_), .A4(new_n384_), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT54), .Z(new_n811_));
  AND2_X1   g610(.A1(new_n413_), .A2(KEYINPUT57), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n374_), .A2(new_n334_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n356_), .A2(new_n375_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n813_), .B(new_n370_), .C1(new_n362_), .C2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n378_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n297_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n383_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n294_), .B1(new_n819_), .B2(new_n381_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n281_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n281_), .B2(new_n823_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n271_), .B(KEYINPUT55), .C1(new_n276_), .C2(new_n280_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n264_), .A2(new_n266_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n270_), .B1(new_n240_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n283_), .B2(KEYINPUT12), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n273_), .B1(new_n829_), .B2(new_n282_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n826_), .A2(new_n830_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n824_), .A2(new_n825_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n821_), .B1(new_n832_), .B2(new_n289_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n826_), .A2(new_n830_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT69), .B1(new_n282_), .B2(new_n273_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n279_), .A2(new_n277_), .A3(new_n272_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n829_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT114), .B1(new_n837_), .B2(KEYINPUT55), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n281_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n834_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n288_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n820_), .B1(new_n833_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n818_), .B1(new_n842_), .B2(KEYINPUT115), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n382_), .A2(new_n383_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n288_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n288_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(KEYINPUT115), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n812_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n294_), .A2(new_n817_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n833_), .B2(new_n841_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT58), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n850_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(KEYINPUT116), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n672_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n818_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n414_), .B1(new_n862_), .B2(new_n847_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n849_), .B(new_n858_), .C1(new_n863_), .C2(KEYINPUT57), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n333_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n809_), .B1(new_n811_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866_), .B2(new_n384_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n810_), .B(KEYINPUT54), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n849_), .A2(new_n858_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n860_), .A2(new_n861_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n847_), .A3(new_n818_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT57), .B1(new_n874_), .B2(new_n413_), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT118), .B(new_n333_), .C1(new_n872_), .C2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n869_), .B1(new_n871_), .B2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n868_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n876_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT118), .B1(new_n864_), .B2(new_n333_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n811_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(KEYINPUT119), .A3(new_n878_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n866_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n880_), .A2(new_n884_), .B1(KEYINPUT59), .B2(new_n885_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n384_), .A2(G113gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n867_), .B1(new_n886_), .B2(new_n887_), .ZN(G1340gat));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n667_), .B1(new_n866_), .B2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n880_), .B2(new_n884_), .ZN(new_n891_));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT120), .B1(new_n892_), .B2(KEYINPUT60), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n304_), .B2(KEYINPUT60), .ZN(new_n894_));
  MUX2_X1   g693(.A(KEYINPUT120), .B(new_n893_), .S(new_n894_), .Z(new_n895_));
  OAI22_X1  g694(.A1(new_n891_), .A2(new_n892_), .B1(new_n885_), .B2(new_n895_), .ZN(G1341gat));
  AOI21_X1  g695(.A(G127gat), .B1(new_n866_), .B2(new_n332_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n332_), .A2(G127gat), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n886_), .B2(new_n898_), .ZN(G1342gat));
  AOI21_X1  g698(.A(G134gat), .B1(new_n866_), .B2(new_n414_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n672_), .A2(G134gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n886_), .B2(new_n901_), .ZN(G1343gat));
  AOI21_X1  g701(.A(new_n658_), .B1(new_n811_), .B2(new_n865_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(new_n680_), .A3(new_n740_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n385_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n509_), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n668_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT121), .B(G148gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1345gat));
  NOR2_X1   g708(.A1(new_n904_), .A2(new_n333_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT61), .B(G155gat), .Z(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1346gat));
  INV_X1    g711(.A(new_n672_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G162gat), .B1(new_n904_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n414_), .A2(new_n519_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n904_), .B2(new_n915_), .ZN(G1347gat));
  INV_X1    g715(.A(KEYINPUT22), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n740_), .A2(new_n680_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n714_), .A2(new_n551_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n883_), .A2(new_n917_), .A3(new_n384_), .A4(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(G169gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n922_), .A2(new_n923_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n922_), .A2(new_n925_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n877_), .A2(new_n385_), .A3(new_n920_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n923_), .B1(new_n928_), .B2(new_n924_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n926_), .B1(new_n927_), .B2(new_n929_), .ZN(G1348gat));
  NOR2_X1   g729(.A1(new_n877_), .A2(new_n920_), .ZN(new_n931_));
  AOI21_X1  g730(.A(G176gat), .B1(new_n931_), .B2(new_n305_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n920_), .B1(new_n811_), .B2(new_n865_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n667_), .A2(G176gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(KEYINPUT123), .B1(new_n933_), .B2(new_n934_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n933_), .A2(KEYINPUT123), .A3(new_n934_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n932_), .A2(new_n935_), .A3(new_n936_), .ZN(G1349gat));
  AOI21_X1  g736(.A(G183gat), .B1(new_n933_), .B2(new_n332_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n333_), .A2(new_n416_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n931_), .B2(new_n939_), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n931_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n877_), .A2(new_n913_), .A3(new_n920_), .ZN(new_n942_));
  INV_X1    g741(.A(G190gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n941_), .B1(new_n942_), .B2(new_n943_), .ZN(G1351gat));
  NAND3_X1  g743(.A1(new_n903_), .A2(new_n384_), .A3(new_n918_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g745(.A(new_n668_), .B1(KEYINPUT124), .B2(G204gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n903_), .A2(new_n918_), .A3(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n949_), .B(KEYINPUT125), .Z(new_n950_));
  XNOR2_X1  g749(.A(new_n948_), .B(new_n950_), .ZN(G1353gat));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952_));
  INV_X1    g751(.A(G211gat), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n332_), .B1(new_n952_), .B2(new_n953_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(KEYINPUT126), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n903_), .A2(new_n918_), .A3(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n952_), .A2(new_n953_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n956_), .B(new_n957_), .ZN(G1354gat));
  INV_X1    g757(.A(G218gat), .ZN(new_n959_));
  NAND4_X1  g758(.A1(new_n903_), .A2(new_n959_), .A3(new_n414_), .A4(new_n918_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n811_), .A2(new_n865_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n658_), .ZN(new_n962_));
  AND4_X1   g761(.A1(new_n672_), .A2(new_n961_), .A3(new_n962_), .A4(new_n918_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n960_), .B1(new_n963_), .B2(new_n959_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(KEYINPUT127), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966_));
  OAI211_X1 g765(.A(new_n966_), .B(new_n960_), .C1(new_n963_), .C2(new_n959_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n967_), .ZN(G1355gat));
endmodule


