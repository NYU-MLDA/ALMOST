//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n583_, new_n584_, new_n585_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT23), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n202_), .B(KEYINPUT79), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(KEYINPUT23), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(G183gat), .B2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  INV_X1    g007(.A(G169gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT80), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(KEYINPUT80), .A3(KEYINPUT22), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n207_), .B(new_n208_), .C1(new_n212_), .C2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n203_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(new_n205_), .B2(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n209_), .A2(new_n216_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(KEYINPUT78), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(KEYINPUT78), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230_));
  INV_X1    g029(.A(G190gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT26), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n231_), .A2(KEYINPUT26), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n229_), .B(new_n232_), .C1(new_n233_), .C2(new_n230_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n227_), .A2(new_n228_), .A3(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n219_), .B1(new_n222_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n236_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT82), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n241_), .B(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G99gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G43gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT31), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n251_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT89), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n258_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n256_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT89), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n255_), .B(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n259_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT90), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT3), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n269_), .A2(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT84), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n270_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT85), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n276_), .B(new_n278_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT83), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(KEYINPUT1), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n281_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n269_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n271_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT29), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G228gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT88), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n268_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n266_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(G228gat), .A3(G233gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n293_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G22gat), .B(G50gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT87), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n288_), .A2(KEYINPUT29), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n288_), .B2(KEYINPUT29), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G78gat), .B(G106gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n299_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n294_), .A2(new_n308_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n300_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n307_), .B1(new_n300_), .B2(new_n309_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n288_), .A2(new_n246_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n245_), .A2(new_n287_), .A3(new_n283_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(KEYINPUT4), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G225gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT94), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n315_), .B(new_n317_), .C1(KEYINPUT4), .C2(new_n313_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n313_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G85gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT0), .B(G57gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  AND3_X1   g122(.A1(new_n318_), .A2(new_n319_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT26), .B(G190gat), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI211_X1 g126(.A(new_n226_), .B(new_n224_), .C1(new_n229_), .C2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n206_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT22), .B(G169gat), .Z(new_n330_));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  OAI221_X1 g130(.A(new_n208_), .B1(G176gat), .B2(new_n330_), .C1(new_n222_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n266_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT20), .B(new_n334_), .C1(new_n268_), .C2(new_n236_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT19), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n268_), .A2(new_n236_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n333_), .A2(new_n266_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n339_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G8gat), .B(G36gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n353_));
  OAI22_X1  g152(.A1(new_n324_), .A2(new_n325_), .B1(new_n346_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n341_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n340_), .A2(KEYINPUT20), .A3(new_n339_), .A4(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n335_), .A2(KEYINPUT92), .A3(new_n337_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT92), .B1(new_n335_), .B2(new_n337_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n353_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT98), .B1(new_n354_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n351_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n352_), .B(new_n356_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n313_), .A2(new_n314_), .A3(new_n317_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n323_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT96), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n315_), .B(new_n316_), .C1(KEYINPUT4), .C2(new_n313_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(KEYINPUT96), .A3(new_n366_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT95), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT33), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n318_), .A2(new_n319_), .A3(new_n323_), .A4(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n318_), .A2(new_n319_), .A3(new_n323_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n363_), .A2(new_n364_), .A3(new_n377_), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n361_), .A2(new_n380_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n354_), .A2(new_n360_), .A3(KEYINPUT98), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n312_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n310_), .A2(new_n311_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n363_), .A2(new_n364_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n324_), .A2(new_n325_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n364_), .B(KEYINPUT27), .C1(new_n352_), .C2(new_n346_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n384_), .A2(new_n387_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n254_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n254_), .A2(new_n388_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n384_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G15gat), .B(G22gat), .ZN(new_n396_));
  INV_X1    g195(.A(G1gat), .ZN(new_n397_));
  INV_X1    g196(.A(G8gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT14), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G8gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G231gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G57gat), .B(G64gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G71gat), .B(G78gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT11), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(KEYINPUT11), .ZN(new_n408_));
  INV_X1    g207(.A(new_n406_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n405_), .A2(KEYINPUT11), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n407_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n404_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G127gat), .B(G155gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT16), .ZN(new_n415_));
  XOR2_X1   g214(.A(G183gat), .B(G211gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n418_));
  OR3_X1    g217(.A1(new_n413_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(KEYINPUT74), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n417_), .B(KEYINPUT17), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n413_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(KEYINPUT74), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G29gat), .B(G36gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G43gat), .B(G50gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT15), .ZN(new_n428_));
  OR2_X1    g227(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n429_));
  INV_X1    g228(.A(G106gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT64), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT64), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n429_), .A2(new_n431_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT65), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT9), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT9), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT65), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n437_), .A2(new_n439_), .A3(G85gat), .A4(G92gat), .ZN(new_n440_));
  INV_X1    g239(.A(G85gat), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n443_), .A2(new_n436_), .A3(KEYINPUT9), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G99gat), .A2(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT6), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(G99gat), .A3(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n435_), .A2(new_n440_), .A3(new_n445_), .A4(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n443_), .A2(new_n444_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI211_X1 g255(.A(KEYINPUT8), .B(new_n452_), .C1(new_n456_), .C2(new_n450_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n430_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n450_), .A2(new_n453_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n452_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n458_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n451_), .B1(new_n457_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n428_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n451_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n447_), .A2(new_n449_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n461_), .A2(new_n453_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n463_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT8), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(new_n458_), .A3(new_n463_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n467_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n427_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n475_));
  NAND2_X1  g274(.A1(G232gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n466_), .A2(new_n474_), .A3(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n477_), .A2(new_n478_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n481_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G190gat), .B(G218gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G134gat), .B(G162gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT36), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n487_), .A2(KEYINPUT36), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n482_), .A2(new_n490_), .A3(new_n483_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n395_), .A2(new_n424_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT69), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT13), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT68), .ZN(new_n497_));
  INV_X1    g296(.A(new_n412_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n465_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n412_), .B(new_n451_), .C1(new_n457_), .C2(new_n464_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(KEYINPUT66), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G230gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n465_), .A2(new_n504_), .A3(new_n498_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n503_), .B1(new_n473_), .B2(new_n412_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n473_), .A2(KEYINPUT12), .A3(new_n412_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT12), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n465_), .B2(new_n498_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n507_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G120gat), .B(G148gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G176gat), .B(G204gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n506_), .A2(new_n511_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n506_), .B2(new_n511_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n497_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n519_), .A2(new_n497_), .A3(new_n520_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n496_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n495_), .A2(KEYINPUT13), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n428_), .A2(new_n402_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT75), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n402_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n533_), .B2(new_n427_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n427_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n402_), .B(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n530_), .A2(new_n534_), .B1(new_n536_), .B2(new_n532_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT76), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G169gat), .B(G197gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n537_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n528_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n494_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(G1gat), .B1(new_n545_), .B2(new_n388_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT100), .Z(new_n547_));
  NOR2_X1   g346(.A1(new_n395_), .A2(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n492_), .A2(KEYINPUT37), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT72), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT71), .B(KEYINPUT37), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n489_), .A2(new_n550_), .A3(new_n491_), .A4(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT72), .B1(new_n492_), .B2(new_n551_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n528_), .A2(new_n556_), .A3(new_n424_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n548_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n388_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n397_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT38), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n547_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT101), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT101), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n547_), .A2(new_n565_), .A3(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(G1324gat));
  NAND3_X1  g366(.A1(new_n559_), .A2(new_n398_), .A3(new_n392_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n545_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n398_), .B1(new_n569_), .B2(new_n392_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT39), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n571_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n568_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n574_), .B(new_n576_), .ZN(G1325gat));
  INV_X1    g376(.A(new_n254_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G15gat), .B1(new_n545_), .B2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT41), .Z(new_n580_));
  NAND3_X1  g379(.A1(new_n559_), .A2(new_n238_), .A3(new_n254_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(G1326gat));
  OAI21_X1  g381(.A(G22gat), .B1(new_n545_), .B2(new_n312_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT42), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n312_), .A2(G22gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n584_), .B1(new_n558_), .B2(new_n585_), .ZN(G1327gat));
  INV_X1    g385(.A(new_n528_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n548_), .A2(new_n587_), .A3(new_n424_), .A4(new_n493_), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n588_), .A2(G29gat), .A3(new_n388_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n424_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n556_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT43), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n556_), .B2(KEYINPUT103), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n590_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n556_), .B(new_n593_), .C1(new_n391_), .C2(new_n394_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n544_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT44), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n595_), .A2(KEYINPUT44), .A3(new_n544_), .A4(new_n596_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n560_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT104), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G29gat), .B1(new_n601_), .B2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n589_), .B1(new_n603_), .B2(new_n604_), .ZN(G1328gat));
  INV_X1    g404(.A(new_n392_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(G36gat), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n588_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT45), .Z(new_n609_));
  NAND3_X1  g408(.A1(new_n599_), .A2(new_n392_), .A3(new_n600_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT105), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G36gat), .B1(new_n610_), .B2(new_n611_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n609_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT46), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n609_), .B(KEYINPUT46), .C1(new_n612_), .C2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1329gat));
  NAND4_X1  g417(.A1(new_n599_), .A2(G43gat), .A3(new_n254_), .A4(new_n600_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT106), .B(G43gat), .Z(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n588_), .B2(new_n578_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g422(.A1(new_n599_), .A2(G50gat), .A3(new_n384_), .A4(new_n600_), .ZN(new_n624_));
  INV_X1    g423(.A(G50gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n588_), .B2(new_n312_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n624_), .A2(new_n626_), .ZN(G1331gat));
  NOR2_X1   g426(.A1(new_n587_), .A2(new_n542_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n494_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G57gat), .B1(new_n629_), .B2(new_n388_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n395_), .A2(new_n542_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n424_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n528_), .A3(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n388_), .A2(G57gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(G1332gat));
  OAI21_X1  g434(.A(G64gat), .B1(new_n629_), .B2(new_n606_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT48), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n606_), .A2(G64gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n633_), .B2(new_n638_), .ZN(G1333gat));
  OAI21_X1  g438(.A(G71gat), .B1(new_n629_), .B2(new_n578_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT49), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n578_), .A2(G71gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n633_), .B2(new_n642_), .ZN(G1334gat));
  OAI21_X1  g442(.A(G78gat), .B1(new_n629_), .B2(new_n312_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT50), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n312_), .A2(G78gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT107), .Z(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n633_), .B2(new_n647_), .ZN(G1335gat));
  NAND4_X1  g447(.A1(new_n631_), .A2(new_n528_), .A3(new_n424_), .A4(new_n493_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n441_), .A3(new_n560_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n595_), .A2(new_n596_), .A3(new_n628_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G85gat), .B1(new_n652_), .B2(new_n388_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1336gat));
  NAND3_X1  g453(.A1(new_n650_), .A2(new_n442_), .A3(new_n392_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G92gat), .B1(new_n652_), .B2(new_n606_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1337gat));
  OAI21_X1  g456(.A(G99gat), .B1(new_n652_), .B2(new_n578_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n254_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n649_), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g460(.A1(new_n650_), .A2(new_n431_), .A3(new_n433_), .A4(new_n384_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n595_), .A2(new_n384_), .A3(new_n596_), .A4(new_n628_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G106gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT108), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT52), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n667_), .A3(G106gat), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n665_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n666_), .B1(new_n665_), .B2(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n662_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT53), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT53), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(new_n662_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1339gat));
  NAND4_X1  g474(.A1(new_n632_), .A2(new_n526_), .A3(new_n543_), .A4(new_n527_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT110), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(KEYINPUT110), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n676_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT57), .ZN(new_n685_));
  INV_X1    g484(.A(new_n523_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n530_), .B(new_n532_), .C1(new_n402_), .C2(new_n535_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n541_), .B1(new_n536_), .B2(new_n531_), .ZN(new_n688_));
  AOI22_X1  g487(.A1(new_n687_), .A2(new_n688_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n686_), .A2(new_n521_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n542_), .A2(new_n518_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT56), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n517_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n500_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n696_));
  AOI22_X1  g495(.A1(new_n503_), .A2(new_n695_), .B1(new_n511_), .B2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT55), .B(new_n507_), .C1(new_n508_), .C2(new_n510_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT112), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(new_n503_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n511_), .A2(new_n696_), .ZN(new_n701_));
  AND4_X1   g500(.A1(KEYINPUT112), .A2(new_n700_), .A3(new_n701_), .A4(new_n698_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n694_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(new_n701_), .A3(new_n698_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n700_), .A2(new_n701_), .A3(new_n698_), .A4(KEYINPUT112), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n517_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n703_), .B1(new_n708_), .B2(KEYINPUT56), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n690_), .B1(new_n692_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n685_), .B1(new_n710_), .B2(new_n493_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n516_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n693_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n691_), .B1(new_n713_), .B2(new_n703_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT57), .B(new_n492_), .C1(new_n714_), .C2(new_n690_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n711_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT113), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n703_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n694_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT113), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n713_), .A2(new_n718_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n689_), .A2(new_n518_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n722_), .A2(KEYINPUT58), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n554_), .A2(new_n555_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(KEYINPUT113), .A2(new_n720_), .B1(new_n708_), .B2(KEYINPUT56), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n703_), .A2(new_n717_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n724_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT58), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n726_), .B1(new_n732_), .B2(KEYINPUT114), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT58), .B1(new_n722_), .B2(new_n724_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n727_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n716_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n684_), .B1(new_n737_), .B2(new_n590_), .ZN(new_n738_));
  NOR4_X1   g537(.A1(new_n392_), .A2(new_n578_), .A3(new_n384_), .A4(new_n388_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(KEYINPUT115), .A3(new_n739_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n542_), .A3(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(G113gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT59), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n717_), .A2(new_n703_), .B1(new_n712_), .B2(new_n693_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n723_), .B1(new_n750_), .B2(new_n721_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT114), .B(new_n556_), .C1(new_n751_), .C2(KEYINPUT58), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n736_), .A2(new_n752_), .A3(new_n725_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n711_), .A2(new_n715_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n590_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n749_), .B(new_n739_), .C1(new_n755_), .C2(new_n683_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n738_), .A2(KEYINPUT117), .A3(new_n749_), .A4(new_n739_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n740_), .A2(KEYINPUT59), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT118), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT118), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n543_), .A2(new_n745_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n748_), .B1(new_n765_), .B2(new_n766_), .ZN(G1340gat));
  INV_X1    g566(.A(KEYINPUT121), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT120), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n587_), .B1(new_n740_), .B2(KEYINPUT59), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n760_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n760_), .B2(new_n770_), .ZN(new_n772_));
  INV_X1    g571(.A(G120gat), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n587_), .A2(KEYINPUT60), .ZN(new_n775_));
  MUX2_X1   g574(.A(KEYINPUT60), .B(new_n775_), .S(new_n773_), .Z(new_n776_));
  NAND3_X1  g575(.A1(new_n742_), .A2(new_n743_), .A3(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT119), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n768_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n777_), .B(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n760_), .A2(new_n770_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G120gat), .B1(new_n782_), .B2(new_n769_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n781_), .B(KEYINPUT121), .C1(new_n783_), .C2(new_n771_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n779_), .A2(new_n784_), .ZN(G1341gat));
  AND2_X1   g584(.A1(new_n742_), .A2(new_n743_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G127gat), .B1(new_n786_), .B2(new_n590_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n424_), .A2(KEYINPUT122), .ZN(new_n788_));
  MUX2_X1   g587(.A(KEYINPUT122), .B(new_n788_), .S(G127gat), .Z(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n765_), .B2(new_n789_), .ZN(G1342gat));
  INV_X1    g589(.A(G134gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n786_), .A2(new_n791_), .A3(new_n493_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n727_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n791_), .ZN(G1343gat));
  INV_X1    g593(.A(new_n738_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n578_), .A2(new_n560_), .A3(new_n384_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n795_), .A2(new_n392_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n542_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n528_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT123), .B(G148gat), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1345gat));
  NAND2_X1  g601(.A1(new_n797_), .A2(new_n590_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(KEYINPUT61), .B(G155gat), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(G1346gat));
  AOI21_X1  g604(.A(G162gat), .B1(new_n797_), .B2(new_n493_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n556_), .A2(G162gat), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT124), .Z(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n797_), .B2(new_n808_), .ZN(G1347gat));
  NOR4_X1   g608(.A1(new_n795_), .A2(new_n384_), .A3(new_n606_), .A4(new_n393_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n209_), .B1(new_n810_), .B2(new_n542_), .ZN(new_n811_));
  XOR2_X1   g610(.A(new_n811_), .B(KEYINPUT62), .Z(new_n812_));
  NOR2_X1   g611(.A1(new_n543_), .A2(new_n330_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT125), .Z(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(G1348gat));
  NAND2_X1  g615(.A1(new_n810_), .A2(new_n528_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g617(.A1(new_n810_), .A2(new_n590_), .ZN(new_n819_));
  MUX2_X1   g618(.A(new_n229_), .B(G183gat), .S(new_n819_), .Z(G1350gat));
  NAND3_X1  g619(.A1(new_n810_), .A2(new_n327_), .A3(new_n493_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n810_), .A2(new_n556_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n821_), .B1(new_n823_), .B2(new_n231_), .ZN(G1351gat));
  NAND3_X1  g623(.A1(new_n578_), .A2(new_n388_), .A3(new_n384_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n392_), .B1(new_n825_), .B2(KEYINPUT126), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n826_), .B(new_n795_), .C1(KEYINPUT126), .C2(new_n825_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n542_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n528_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n590_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n833_));
  AND2_X1   g632(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n832_), .B2(new_n833_), .ZN(G1354gat));
  NAND2_X1  g635(.A1(new_n827_), .A2(new_n493_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT127), .B(G218gat), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n727_), .A2(new_n838_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n837_), .A2(new_n838_), .B1(new_n827_), .B2(new_n839_), .ZN(G1355gat));
endmodule


