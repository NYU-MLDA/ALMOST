//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT89), .B(G204gat), .Z(new_n203_));
  INV_X1    g002(.A(G197gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT90), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT90), .ZN(new_n208_));
  NOR3_X1   g007(.A1(new_n203_), .A2(new_n208_), .A3(G197gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(KEYINPUT21), .B(new_n202_), .C1(new_n207_), .C2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT91), .A2(KEYINPUT21), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n202_), .B(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n204_), .A2(G204gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n203_), .A2(G197gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  INV_X1    g018(.A(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT81), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  OR3_X1    g023(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT22), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT22), .B1(new_n223_), .B2(new_n224_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n222_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT24), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(KEYINPUT24), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(new_n231_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(KEYINPUT80), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT26), .B(G190gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT80), .B1(new_n219_), .B2(KEYINPUT25), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n218_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n230_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n216_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n222_), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT22), .B(G169gat), .Z(new_n245_));
  OAI21_X1  g044(.A(new_n229_), .B1(new_n245_), .B2(G176gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n236_), .A2(new_n238_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n218_), .ZN(new_n248_));
  OAI22_X1  g047(.A1(new_n244_), .A2(new_n246_), .B1(new_n248_), .B2(new_n235_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n243_), .B(KEYINPUT20), .C1(new_n216_), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G226gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT19), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n216_), .A2(new_n249_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n254_), .B(KEYINPUT20), .C1(new_n242_), .C2(new_n216_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G8gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT94), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G64gat), .B(G92gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT95), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT95), .B1(new_n256_), .B2(new_n262_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G225gat), .A2(G233gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(G155gat), .B2(G162gat), .ZN(new_n273_));
  OR2_X1    g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT85), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(KEYINPUT3), .Z(new_n276_));
  NAND2_X1  g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT2), .Z(new_n278_));
  OAI21_X1  g077(.A(new_n273_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(G155gat), .B2(G162gat), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n272_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(G155gat), .A3(G162gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT84), .Z(new_n284_));
  OAI211_X1 g083(.A(new_n277_), .B(new_n274_), .C1(new_n282_), .C2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G127gat), .B(G134gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n286_), .A2(KEYINPUT4), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n286_), .B(new_n289_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT4), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n269_), .B(new_n290_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n279_), .A2(new_n285_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(new_n289_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n268_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G29gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT0), .ZN(new_n298_));
  INV_X1    g097(.A(G57gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G85gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n293_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT33), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n304_), .A2(new_n305_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n291_), .A2(new_n292_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n290_), .A2(new_n268_), .ZN(new_n309_));
  OAI221_X1 g108(.A(new_n302_), .B1(new_n291_), .B2(new_n268_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n267_), .A2(new_n306_), .A3(new_n307_), .A4(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n293_), .A2(new_n296_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n302_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n313_), .A2(new_n304_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n250_), .A2(KEYINPUT96), .A3(new_n252_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT96), .B1(new_n250_), .B2(new_n252_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(KEYINPUT32), .A3(new_n262_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n262_), .A2(KEYINPUT32), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n256_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n311_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n216_), .B1(new_n286_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327_));
  OR2_X1    g126(.A1(KEYINPUT88), .A2(G228gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(KEYINPUT88), .A2(G228gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n216_), .A2(new_n327_), .B1(G233gat), .B2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n326_), .B(new_n331_), .Z(new_n332_));
  XNOR2_X1  g131(.A(G78gat), .B(G106gat), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n334_), .A2(KEYINPUT93), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n326_), .B(new_n331_), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n333_), .B(KEYINPUT92), .Z(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n294_), .A2(KEYINPUT29), .ZN(new_n339_));
  XOR2_X1   g138(.A(G22gat), .B(G50gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n334_), .A2(KEYINPUT93), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n335_), .A2(new_n338_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n336_), .B(new_n337_), .Z(new_n346_));
  OR2_X1    g145(.A1(new_n346_), .A2(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT97), .B1(new_n324_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n323_), .B2(new_n311_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT97), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n267_), .A2(KEYINPUT27), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n319_), .A2(new_n261_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(KEYINPUT27), .A3(new_n263_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(new_n314_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n349_), .B(new_n352_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G43gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G15gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n361_), .B(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n359_), .B(new_n365_), .Z(new_n366_));
  XOR2_X1   g165(.A(new_n289_), .B(KEYINPUT31), .Z(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(KEYINPUT82), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n366_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n356_), .A2(new_n348_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n315_), .A2(new_n370_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n358_), .A2(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G141gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT79), .ZN(new_n375_));
  XOR2_X1   g174(.A(G169gat), .B(G197gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G29gat), .B(G36gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n378_), .A2(new_n379_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G43gat), .B(G50gat), .Z(new_n382_));
  OR3_X1    g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT15), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G1gat), .B(G8gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT78), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G15gat), .B(G22gat), .ZN(new_n390_));
  INV_X1    g189(.A(G1gat), .ZN(new_n391_));
  INV_X1    g190(.A(G8gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT14), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n389_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n387_), .A2(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n395_), .A2(new_n385_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G229gat), .A2(G233gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n383_), .A2(new_n384_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(new_n395_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n377_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n404_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n377_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT7), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT7), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT65), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G99gat), .A2(G106gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n412_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n413_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G99gat), .A2(G106gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT6), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(G99gat), .A3(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT8), .ZN(new_n425_));
  XOR2_X1   g224(.A(G85gat), .B(G92gat), .Z(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(KEYINPUT66), .A2(KEYINPUT67), .ZN(new_n428_));
  NOR2_X1   g227(.A1(KEYINPUT66), .A2(KEYINPUT67), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n420_), .B(new_n422_), .C1(new_n429_), .C2(new_n428_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n418_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT68), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n426_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT8), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n434_), .B1(new_n433_), .B2(new_n426_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n427_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G57gat), .B(G64gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT11), .ZN(new_n440_));
  XOR2_X1   g239(.A(G71gat), .B(G78gat), .Z(new_n441_));
  OR2_X1    g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n441_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n439_), .A2(KEYINPUT11), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT10), .B(G99gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT64), .ZN(new_n447_));
  INV_X1    g246(.A(G106gat), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n426_), .A2(KEYINPUT9), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G85gat), .A2(G92gat), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n450_), .B(new_n423_), .C1(KEYINPUT9), .C2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n438_), .A2(new_n445_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT69), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n433_), .A2(new_n426_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT68), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(KEYINPUT8), .A3(new_n435_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n453_), .B1(new_n460_), .B2(new_n427_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT69), .A3(new_n445_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n438_), .A2(new_n454_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n445_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n457_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(G230gat), .A2(G233gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n461_), .B2(new_n445_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n467_), .B1(new_n461_), .B2(new_n445_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n438_), .A2(KEYINPUT70), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT70), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(new_n427_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n453_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n464_), .A2(KEYINPUT12), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n470_), .B(new_n471_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G120gat), .B(G148gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT5), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G176gat), .B(G204gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n468_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT72), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n468_), .A2(KEYINPUT72), .A3(new_n477_), .A4(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n468_), .A2(new_n477_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n487_), .B1(new_n488_), .B2(new_n482_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT73), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT35), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G232gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT34), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n461_), .A2(new_n401_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n387_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(new_n475_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n496_), .A2(new_n493_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G190gat), .B(G218gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT75), .ZN(new_n503_));
  XOR2_X1   g302(.A(G134gat), .B(G162gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n500_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n497_), .B(new_n508_), .C1(new_n475_), .C2(new_n498_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n501_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT76), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n501_), .A2(new_n512_), .A3(new_n507_), .A4(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n505_), .B(new_n506_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n501_), .B2(new_n509_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT37), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n514_), .A2(new_n517_), .A3(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G231gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n395_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(new_n464_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529_));
  XOR2_X1   g328(.A(G127gat), .B(G155gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT16), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G183gat), .B(G211gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n528_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(KEYINPUT17), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n524_), .A2(new_n538_), .ZN(new_n539_));
  NOR4_X1   g338(.A1(new_n373_), .A2(new_n410_), .A3(new_n492_), .A4(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n391_), .A3(new_n315_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT38), .ZN(new_n542_));
  OAI22_X1  g341(.A1(new_n350_), .A2(new_n351_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n324_), .A2(KEYINPUT97), .A3(new_n348_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n370_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n371_), .A2(new_n372_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n491_), .A2(new_n410_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n537_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(G1gat), .B1(new_n552_), .B2(new_n314_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n542_), .A2(new_n553_), .ZN(G1324gat));
  AOI21_X1  g353(.A(new_n392_), .B1(new_n551_), .B2(new_n356_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT39), .Z(new_n556_));
  NAND3_X1  g355(.A1(new_n540_), .A2(new_n392_), .A3(new_n356_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT40), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(KEYINPUT40), .A3(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(G1325gat));
  OAI21_X1  g361(.A(G15gat), .B1(new_n552_), .B2(new_n370_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT41), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(KEYINPUT41), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n540_), .A2(new_n363_), .A3(new_n369_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(G1326gat));
  INV_X1    g366(.A(G22gat), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n551_), .B2(new_n348_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT42), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n348_), .A2(new_n568_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT98), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n540_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(G1327gat));
  NOR2_X1   g373(.A1(new_n518_), .A2(new_n538_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n549_), .A2(KEYINPUT101), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n547_), .A2(new_n548_), .A3(new_n575_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(G29gat), .B1(new_n581_), .B2(new_n315_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n548_), .A2(new_n537_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT99), .Z(new_n584_));
  INV_X1    g383(.A(KEYINPUT43), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n514_), .A2(new_n517_), .A3(new_n520_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n520_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n585_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n373_), .B2(new_n524_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n547_), .B(new_n588_), .C1(new_n589_), .C2(new_n585_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n584_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT44), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(KEYINPUT44), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n596_), .A2(G29gat), .A3(new_n315_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n582_), .B1(new_n595_), .B2(new_n597_), .ZN(G1328gat));
  INV_X1    g397(.A(new_n356_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(G36gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n576_), .A2(new_n579_), .A3(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT45), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(KEYINPUT45), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n596_), .A2(new_n356_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G36gat), .B1(new_n605_), .B2(new_n594_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n604_), .B(new_n606_), .C1(KEYINPUT102), .C2(KEYINPUT46), .ZN(new_n607_));
  NAND2_X1  g406(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(G1329gat));
  NAND3_X1  g408(.A1(new_n596_), .A2(G43gat), .A3(new_n369_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n580_), .A2(new_n370_), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n610_), .A2(new_n594_), .B1(new_n611_), .B2(G43gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT103), .B(KEYINPUT47), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(G1330gat));
  NAND2_X1  g413(.A1(new_n596_), .A2(new_n348_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G50gat), .B1(new_n615_), .B2(new_n594_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n348_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(G50gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT104), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n616_), .B1(new_n580_), .B2(new_n619_), .ZN(G1331gat));
  AND2_X1   g419(.A1(new_n491_), .A2(new_n410_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n547_), .A2(new_n538_), .A3(new_n524_), .A4(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT105), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n299_), .A3(new_n315_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n410_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n492_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n373_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n550_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G57gat), .B1(new_n628_), .B2(new_n314_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n624_), .A2(new_n629_), .ZN(G1332gat));
  OAI21_X1  g429(.A(G64gat), .B1(new_n628_), .B2(new_n599_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT48), .ZN(new_n632_));
  INV_X1    g431(.A(G64gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n623_), .A2(new_n633_), .A3(new_n356_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1333gat));
  OAI21_X1  g434(.A(G71gat), .B1(new_n628_), .B2(new_n370_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT49), .ZN(new_n637_));
  INV_X1    g436(.A(G71gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n623_), .A2(new_n638_), .A3(new_n369_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1334gat));
  OAI21_X1  g439(.A(G78gat), .B1(new_n628_), .B2(new_n617_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT50), .ZN(new_n642_));
  INV_X1    g441(.A(G78gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n623_), .A2(new_n643_), .A3(new_n348_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1335gat));
  NAND2_X1  g444(.A1(new_n627_), .A2(new_n575_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G85gat), .B1(new_n647_), .B2(new_n315_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n621_), .A2(new_n537_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n315_), .A2(G85gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT106), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n648_), .B1(new_n650_), .B2(new_n652_), .ZN(G1336gat));
  AOI21_X1  g452(.A(G92gat), .B1(new_n647_), .B2(new_n356_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT107), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n356_), .A2(G92gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT108), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n650_), .B2(new_n657_), .ZN(G1337gat));
  INV_X1    g457(.A(KEYINPUT110), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n650_), .A2(new_n369_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n369_), .A2(new_n447_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n660_), .A2(G99gat), .B1(new_n647_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT109), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n662_), .A2(KEYINPUT109), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n659_), .B(KEYINPUT51), .C1(new_n664_), .C2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT51), .ZN(new_n667_));
  INV_X1    g466(.A(new_n665_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(new_n663_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT110), .B1(new_n662_), .B2(new_n667_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(G1338gat));
  NAND3_X1  g470(.A1(new_n647_), .A2(new_n448_), .A3(new_n348_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT52), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n650_), .A2(new_n674_), .A3(new_n348_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G106gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n674_), .B1(new_n650_), .B2(new_n348_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n673_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n676_), .A2(KEYINPUT52), .A3(new_n678_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n672_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT53), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT53), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(new_n672_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1339gat));
  NOR3_X1   g485(.A1(new_n539_), .A2(new_n491_), .A3(new_n625_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT54), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n398_), .A2(new_n399_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n377_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(new_n691_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n405_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n489_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n470_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n457_), .A2(new_n462_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n467_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n474_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n473_), .B1(new_n460_), .B2(new_n427_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n454_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n476_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n704_), .A2(KEYINPUT55), .A3(new_n470_), .A4(new_n471_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT55), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n477_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n699_), .A2(new_n705_), .A3(new_n707_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n708_), .A2(KEYINPUT56), .A3(new_n481_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT56), .B1(new_n708_), .B2(new_n481_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n410_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n709_), .A2(new_n710_), .B1(new_n711_), .B2(KEYINPUT112), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(KEYINPUT112), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n696_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n518_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT57), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT58), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n709_), .A2(new_n710_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n487_), .A2(new_n695_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT114), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n588_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n708_), .A2(new_n481_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT56), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n708_), .A2(KEYINPUT56), .A3(new_n481_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n487_), .A2(new_n695_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(KEYINPUT58), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n723_), .A2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n722_), .B1(new_n721_), .B2(new_n588_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n717_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT116), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n715_), .A2(new_n716_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT58), .B1(new_n728_), .B2(new_n729_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT114), .B1(new_n524_), .B2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n723_), .A3(new_n730_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(KEYINPUT116), .A3(new_n717_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n735_), .A2(new_n737_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n537_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(new_n537_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n689_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n371_), .A2(new_n315_), .A3(new_n369_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(KEYINPUT59), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n537_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n689_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n747_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT59), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n749_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G113gat), .B1(new_n755_), .B2(new_n410_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n753_), .B(KEYINPUT115), .Z(new_n757_));
  INV_X1    g556(.A(G113gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n625_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(G1340gat));
  AND3_X1   g559(.A1(new_n740_), .A2(KEYINPUT116), .A3(new_n717_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT116), .B1(new_n740_), .B2(new_n717_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n736_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT117), .B1(new_n763_), .B2(new_n538_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n742_), .A2(new_n743_), .A3(new_n537_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n688_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n748_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n492_), .B(new_n754_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n749_), .A2(KEYINPUT118), .A3(new_n492_), .A4(new_n754_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(G120gat), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT60), .ZN(new_n773_));
  INV_X1    g572(.A(G120gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n491_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n757_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n772_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT119), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n772_), .A2(new_n780_), .A3(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1341gat));
  AOI21_X1  g581(.A(G127gat), .B1(new_n757_), .B2(new_n538_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n755_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n538_), .A2(G127gat), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT120), .Z(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n784_), .B2(new_n786_), .ZN(G1342gat));
  INV_X1    g586(.A(G134gat), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n757_), .A2(new_n788_), .A3(new_n514_), .A4(new_n517_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n755_), .A2(new_n524_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(new_n788_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT121), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n789_), .B(KEYINPUT121), .C1(new_n790_), .C2(new_n788_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1343gat));
  AOI211_X1 g594(.A(new_n369_), .B(new_n617_), .C1(new_n689_), .C2(new_n750_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n356_), .A2(new_n314_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n625_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n492_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n538_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT122), .ZN(new_n805_));
  XOR2_X1   g604(.A(KEYINPUT61), .B(G155gat), .Z(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1346gat));
  OAI21_X1  g606(.A(G162gat), .B1(new_n798_), .B2(new_n524_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n518_), .A2(G162gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n798_), .B2(new_n809_), .ZN(G1347gat));
  NAND2_X1  g609(.A1(new_n746_), .A2(new_n617_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n356_), .A2(new_n372_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n625_), .ZN(new_n814_));
  OR3_X1    g613(.A1(new_n811_), .A2(new_n245_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n814_), .B(KEYINPUT123), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n746_), .A2(new_n816_), .A3(new_n617_), .A4(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(G169gat), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT124), .B1(new_n811_), .B2(new_n817_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n815_), .B1(new_n823_), .B2(new_n824_), .ZN(G1348gat));
  NOR2_X1   g624(.A1(new_n811_), .A2(new_n812_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G176gat), .B1(new_n826_), .B2(new_n491_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n751_), .A2(new_n617_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n626_), .A2(new_n226_), .A3(new_n812_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n827_), .B1(new_n829_), .B2(new_n830_), .ZN(G1349gat));
  NOR2_X1   g630(.A1(new_n537_), .A2(new_n236_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n538_), .A3(new_n813_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n826_), .A2(new_n832_), .B1(new_n219_), .B2(new_n833_), .ZN(G1350gat));
  NAND3_X1  g633(.A1(new_n514_), .A2(new_n517_), .A3(new_n238_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT125), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n826_), .A2(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n811_), .A2(new_n524_), .A3(new_n812_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n220_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT126), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT126), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n837_), .B(new_n841_), .C1(new_n220_), .C2(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1351gat));
  NAND3_X1  g642(.A1(new_n796_), .A2(new_n314_), .A3(new_n356_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n410_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(new_n204_), .ZN(G1352gat));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n626_), .ZN(new_n847_));
  MUX2_X1   g646(.A(G204gat), .B(new_n203_), .S(new_n847_), .Z(G1353gat));
  NOR2_X1   g647(.A1(new_n844_), .A2(new_n537_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n850_));
  AND2_X1   g649(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n849_), .B2(new_n850_), .ZN(G1354gat));
  INV_X1    g652(.A(G218gat), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n844_), .A2(new_n854_), .A3(new_n524_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n844_), .A2(new_n518_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n856_), .A2(KEYINPUT127), .ZN(new_n857_));
  AOI21_X1  g656(.A(G218gat), .B1(new_n856_), .B2(KEYINPUT127), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n855_), .B1(new_n857_), .B2(new_n858_), .ZN(G1355gat));
endmodule


