//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G155gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT16), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G211gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT17), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G15gat), .B(G22gat), .Z(new_n210_));
  NAND2_X1  g009(.A1(G1gat), .A2(G8gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(KEYINPUT14), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT72), .ZN(new_n213_));
  XOR2_X1   g012(.A(G1gat), .B(G8gat), .Z(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G57gat), .B(G64gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT11), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G71gat), .B(G78gat), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n216_), .A2(KEYINPUT11), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n218_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n215_), .B(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n209_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n207_), .A2(new_n208_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT37), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT10), .B(G99gat), .Z(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G85gat), .B(G92gat), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT9), .ZN(new_n237_));
  INV_X1    g036(.A(G85gat), .ZN(new_n238_));
  INV_X1    g037(.A(G92gat), .ZN(new_n239_));
  OR3_X1    g038(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT9), .ZN(new_n240_));
  AND3_X1   g039(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n235_), .A2(new_n237_), .A3(new_n240_), .A4(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G99gat), .A2(G106gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(KEYINPUT65), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(new_n252_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n236_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n246_), .B1(new_n259_), .B2(KEYINPUT8), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT8), .ZN(new_n261_));
  AOI211_X1 g060(.A(KEYINPUT66), .B(new_n261_), .C1(new_n258_), .C2(new_n236_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n250_), .A2(new_n243_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(new_n261_), .A3(new_n236_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n245_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G29gat), .ZN(new_n267_));
  INV_X1    g066(.A(G36gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G43gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G29gat), .A2(G36gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G50gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n270_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n269_), .A2(new_n271_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G43gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(G50gat), .B1(new_n278_), .B2(new_n272_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n266_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n259_), .A2(KEYINPUT8), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT66), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n259_), .A2(new_n246_), .A3(KEYINPUT8), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n265_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n244_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n274_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n278_), .A2(G50gat), .A3(new_n272_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n288_), .A2(KEYINPUT15), .A3(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT15), .B1(new_n288_), .B2(new_n289_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n282_), .B1(new_n287_), .B2(new_n293_), .ZN(new_n294_));
  AOI211_X1 g093(.A(KEYINPUT69), .B(new_n292_), .C1(new_n286_), .C2(new_n244_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n281_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G232gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT34), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(KEYINPUT35), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT69), .B1(new_n266_), .B2(new_n292_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n287_), .A2(new_n282_), .A3(new_n293_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n298_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT35), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n304_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n302_), .A2(new_n306_), .A3(new_n307_), .A4(new_n281_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n299_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G190gat), .B(G218gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(G134gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G162gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT36), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT71), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(KEYINPUT71), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n309_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n312_), .A2(KEYINPUT36), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT70), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n299_), .A2(new_n308_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n232_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n299_), .A2(new_n308_), .A3(new_n320_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n314_), .B1(new_n299_), .B2(new_n308_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n323_), .A2(new_n324_), .A3(KEYINPUT37), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n231_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT74), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n231_), .B(new_n328_), .C1(new_n322_), .C2(new_n325_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT13), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G176gat), .B(G204gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G120gat), .B(G148gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G230gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT64), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n265_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n260_), .A2(new_n262_), .A3(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n222_), .B1(new_n341_), .B2(new_n245_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n222_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n286_), .A2(new_n244_), .A3(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(KEYINPUT12), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT12), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n287_), .A2(new_n346_), .A3(new_n222_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n339_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n338_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n336_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n348_), .A2(new_n349_), .A3(new_n336_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n330_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OR3_X1    g152(.A1(new_n348_), .A2(new_n349_), .A3(new_n336_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(KEYINPUT13), .A3(new_n350_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n353_), .A2(KEYINPUT68), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT68), .B1(new_n353_), .B2(new_n355_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n327_), .A2(KEYINPUT75), .A3(new_n329_), .A4(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n213_), .A2(new_n214_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n213_), .A2(new_n214_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n280_), .B(KEYINPUT76), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n215_), .A2(new_n363_), .ZN(new_n366_));
  OAI211_X1 g165(.A(G229gat), .B(G233gat), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n215_), .A2(new_n293_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G229gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT77), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G113gat), .B(G141gat), .ZN(new_n375_));
  INV_X1    g174(.A(G169gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G197gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n367_), .A2(new_n373_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n359_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G1gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(G78gat), .B(G106gat), .Z(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(G228gat), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT89), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(G155gat), .B2(G162gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(KEYINPUT82), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT1), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT83), .ZN(new_n399_));
  OR3_X1    g198(.A1(new_n395_), .A2(new_n397_), .A3(KEYINPUT1), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(KEYINPUT1), .C1(new_n395_), .C2(new_n397_), .ZN(new_n402_));
  OR2_X1    g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n399_), .A2(new_n400_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G141gat), .ZN(new_n405_));
  INV_X1    g204(.A(G148gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT84), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT84), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(G141gat), .B2(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n410_), .A2(new_n412_), .A3(KEYINPUT85), .A4(new_n413_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n407_), .A2(KEYINPUT3), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n408_), .B(KEYINPUT2), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .A4(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n403_), .C1(new_n395_), .C2(new_n397_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n409_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT29), .ZN(new_n423_));
  XOR2_X1   g222(.A(G197gat), .B(G204gat), .Z(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT21), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G197gat), .B(G204gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT21), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G211gat), .B(G218gat), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n425_), .A2(KEYINPUT88), .A3(new_n428_), .A4(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(KEYINPUT88), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(KEYINPUT21), .A3(new_n424_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n393_), .B1(new_n423_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n409_), .B2(new_n421_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n433_), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n391_), .B(KEYINPUT89), .Z(new_n438_));
  NOR3_X1   g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n387_), .B1(new_n434_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n441_));
  INV_X1    g240(.A(new_n438_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n423_), .A2(new_n433_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n392_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n386_), .A3(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G22gat), .B(G50gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n422_), .B2(KEYINPUT29), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n409_), .A2(new_n421_), .A3(new_n435_), .A4(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n447_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(KEYINPUT90), .B(new_n387_), .C1(new_n434_), .C2(new_n439_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n446_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n440_), .A2(new_n445_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT91), .B1(new_n458_), .B2(new_n455_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n454_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(new_n452_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n445_), .A4(new_n440_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n459_), .A3(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G71gat), .B(G99gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT30), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G227gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G15gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n466_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G183gat), .A2(G190gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT23), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT78), .B(G183gat), .Z(new_n473_));
  OAI21_X1  g272(.A(new_n472_), .B1(G190gat), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT79), .ZN(new_n475_));
  OR3_X1    g274(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT79), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n472_), .B(new_n477_), .C1(G190gat), .C2(new_n473_), .ZN(new_n478_));
  OAI21_X1  g277(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n475_), .A2(new_n476_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT26), .B(G190gat), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n473_), .A2(KEYINPUT25), .ZN(new_n482_));
  NOR2_X1   g281(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G176gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n376_), .A2(new_n485_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n486_), .A2(KEYINPUT24), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G169gat), .A2(G176gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(KEYINPUT24), .A3(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n472_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n484_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n480_), .A2(new_n491_), .A3(new_n270_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n270_), .B1(new_n480_), .B2(new_n491_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n470_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n494_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n492_), .A3(new_n469_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT81), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n497_), .A3(KEYINPUT81), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G127gat), .B(G134gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G113gat), .B(G120gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT80), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n502_), .A2(new_n503_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n506_), .A2(KEYINPUT80), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT31), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n500_), .A2(new_n501_), .A3(new_n509_), .ZN(new_n510_));
  OR3_X1    g309(.A1(new_n498_), .A2(new_n499_), .A3(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n464_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n510_), .A2(new_n511_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n514_), .A2(new_n457_), .A3(new_n459_), .A4(new_n463_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n409_), .A2(new_n504_), .A3(new_n421_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n508_), .B1(new_n409_), .B2(new_n421_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n508_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n422_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G225gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n516_), .B1(new_n520_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n422_), .A2(new_n521_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n504_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n527_), .B(KEYINPUT4), .C1(new_n528_), .C2(new_n422_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n523_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(KEYINPUT94), .A3(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n517_), .A2(new_n518_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n523_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n526_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n535_));
  XNOR2_X1  g334(.A(G1gat), .B(G29gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G85gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  OR3_X1    g338(.A1(new_n534_), .A2(KEYINPUT98), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(new_n539_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n539_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n526_), .A2(new_n531_), .A3(new_n542_), .A4(new_n533_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(KEYINPUT98), .A3(new_n543_), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n513_), .A2(new_n515_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G226gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT19), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n472_), .B1(G183gat), .B2(G190gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT22), .B(G169gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT92), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n488_), .B(new_n549_), .C1(new_n551_), .C2(G176gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT25), .B(G183gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n481_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n490_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n548_), .B1(new_n556_), .B2(new_n437_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT96), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n480_), .A2(new_n491_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n433_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n547_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n552_), .A2(new_n555_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n433_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n437_), .A2(new_n480_), .A3(new_n491_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n547_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(KEYINPUT20), .A4(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT97), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(KEYINPUT97), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G8gat), .B(G36gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT18), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G64gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n239_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n557_), .A2(new_n567_), .A3(new_n561_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n565_), .A2(new_n566_), .A3(KEYINPUT20), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n547_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n580_), .A3(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(KEYINPUT27), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n580_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n576_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(KEYINPUT93), .A3(new_n581_), .ZN(new_n585_));
  OR3_X1    g384(.A1(new_n583_), .A2(KEYINPUT93), .A3(new_n576_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT27), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n575_), .A2(KEYINPUT32), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n583_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n571_), .B2(new_n590_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n544_), .A2(new_n540_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n543_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n529_), .A2(new_n523_), .A3(new_n522_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n532_), .A2(new_n524_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n539_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n585_), .A2(new_n586_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n543_), .A2(new_n594_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(new_n598_), .A3(new_n599_), .A4(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n464_), .A2(new_n514_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n545_), .A2(new_n589_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n327_), .A2(new_n329_), .A3(new_n358_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n544_), .A2(new_n540_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n384_), .A2(new_n385_), .A3(new_n607_), .A4(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT99), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n610_), .A2(KEYINPUT99), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n202_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(KEYINPUT38), .A3(new_n611_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n353_), .A2(new_n355_), .A3(new_n383_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT100), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n323_), .A2(new_n324_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n353_), .A2(new_n620_), .A3(new_n355_), .A4(new_n383_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n513_), .A2(new_n515_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n608_), .A3(new_n589_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n602_), .A2(new_n603_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n229_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n608_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT101), .Z(new_n630_));
  NAND3_X1  g429(.A1(new_n614_), .A2(new_n616_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT102), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n614_), .A2(new_n616_), .A3(new_n633_), .A4(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1324gat));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n605_), .A2(new_n606_), .ZN(new_n638_));
  AND4_X1   g437(.A1(new_n638_), .A2(new_n626_), .A3(new_n359_), .A4(new_n383_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640_));
  INV_X1    g439(.A(G8gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n589_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .A4(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n384_), .A2(new_n641_), .A3(new_n607_), .A4(new_n642_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT103), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n622_), .A2(new_n626_), .A3(new_n627_), .A4(new_n642_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(G8gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G8gat), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n637_), .B1(new_n646_), .B2(new_n652_), .ZN(new_n653_));
  AOI211_X1 g452(.A(KEYINPUT104), .B(new_n651_), .C1(new_n643_), .C2(new_n645_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n636_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n644_), .A2(KEYINPUT103), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n644_), .A2(KEYINPUT103), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n652_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT104), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n646_), .A2(new_n637_), .A3(new_n652_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(KEYINPUT40), .A3(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n655_), .A2(new_n661_), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n628_), .B2(new_n512_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT41), .Z(new_n664_));
  INV_X1    g463(.A(new_n639_), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n665_), .A2(G15gat), .A3(new_n512_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(KEYINPUT105), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(KEYINPUT105), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(G1326gat));
  INV_X1    g468(.A(new_n464_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G22gat), .B1(new_n628_), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT42), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n670_), .A2(G22gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n665_), .B2(new_n673_), .ZN(G1327gat));
  NOR2_X1   g473(.A1(new_n604_), .A2(new_n617_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n231_), .A2(new_n619_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n267_), .A3(new_n609_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n323_), .A2(new_n324_), .A3(KEYINPUT37), .ZN(new_n680_));
  INV_X1    g479(.A(new_n315_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n681_), .B(new_n316_), .C1(new_n299_), .C2(new_n308_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT37), .B1(new_n682_), .B2(new_n323_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n679_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n604_), .C2(new_n684_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n231_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n618_), .A2(new_n691_), .A3(new_n621_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT106), .Z(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n690_), .A2(new_n693_), .A3(new_n695_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n608_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n678_), .B1(new_n699_), .B2(new_n267_), .ZN(G1328gat));
  XOR2_X1   g499(.A(new_n589_), .B(KEYINPUT109), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n677_), .A2(new_n268_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT110), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n677_), .A2(new_n704_), .A3(new_n268_), .A4(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n589_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n707_), .B(KEYINPUT46), .C1(new_n268_), .C2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n706_), .B(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n708_), .A2(new_n268_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n709_), .A2(new_n714_), .ZN(G1329gat));
  XOR2_X1   g514(.A(KEYINPUT112), .B(G43gat), .Z(new_n716_));
  INV_X1    g515(.A(new_n677_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n512_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n697_), .A2(new_n698_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n512_), .A2(new_n270_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT111), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n690_), .A2(new_n695_), .A3(new_n693_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n695_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT111), .B(new_n720_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n718_), .B1(new_n721_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT47), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n728_), .B(new_n718_), .C1(new_n721_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1330gat));
  NAND3_X1  g529(.A1(new_n677_), .A2(new_n274_), .A3(new_n464_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n670_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n274_), .ZN(G1331gat));
  NOR2_X1   g532(.A1(new_n358_), .A2(new_n383_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n626_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n619_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n691_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n608_), .B2(KEYINPUT113), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n737_), .B(new_n738_), .C1(KEYINPUT113), .C2(G57gat), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n353_), .A2(new_n355_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n383_), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n327_), .A2(new_n626_), .A3(new_n329_), .A4(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n608_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n739_), .B1(new_n744_), .B2(G57gat), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT114), .ZN(G1332gat));
  INV_X1    g545(.A(new_n737_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n701_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G64gat), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT48), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(G64gat), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT115), .Z(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n743_), .B2(new_n752_), .ZN(G1333gat));
  OR3_X1    g552(.A1(new_n743_), .A2(G71gat), .A3(new_n512_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G71gat), .B1(new_n747_), .B2(new_n512_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n755_), .A2(KEYINPUT116), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(KEYINPUT116), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(KEYINPUT49), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT49), .B1(new_n756_), .B2(new_n757_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n758_), .B2(new_n759_), .ZN(G1334gat));
  OAI21_X1  g559(.A(G78gat), .B1(new_n747_), .B2(new_n670_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT50), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n670_), .A2(G78gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n743_), .B2(new_n763_), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n735_), .A2(new_n619_), .A3(new_n231_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n609_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n690_), .A2(new_n691_), .A3(new_n741_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n608_), .A2(new_n238_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(G1336gat));
  AOI21_X1  g568(.A(G92gat), .B1(new_n765_), .B2(new_n642_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n748_), .A2(new_n239_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n767_), .B2(new_n771_), .ZN(G1337gat));
  NAND2_X1  g571(.A1(new_n767_), .A2(new_n514_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G99gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n765_), .A2(new_n233_), .A3(new_n514_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT117), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n776_), .B(new_n778_), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n234_), .A3(new_n464_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n690_), .A2(new_n691_), .A3(new_n464_), .A4(new_n741_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g585(.A1(new_n642_), .A2(new_n515_), .A3(new_n608_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n372_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n368_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n379_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT118), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n789_), .A2(new_n793_), .A3(new_n379_), .A4(new_n790_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n382_), .A3(new_n794_), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n795_), .A2(KEYINPUT119), .A3(new_n352_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT119), .B1(new_n795_), .B2(new_n352_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n348_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n799_), .A2(KEYINPUT55), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n345_), .A2(new_n339_), .A3(new_n347_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(KEYINPUT55), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n336_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n336_), .A4(new_n802_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n803_), .A2(KEYINPUT120), .A3(new_n804_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n798_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n684_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n798_), .A2(new_n808_), .A3(KEYINPUT58), .A4(new_n809_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n383_), .A2(new_n354_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n795_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n619_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n619_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n815_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n229_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n383_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n684_), .A2(new_n231_), .A3(new_n740_), .A4(new_n826_), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT54), .Z(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n788_), .B1(new_n825_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830_), .B2(new_n383_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n231_), .B1(new_n815_), .B2(new_n823_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(new_n828_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n788_), .A2(KEYINPUT59), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n627_), .B1(new_n815_), .B2(new_n823_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n787_), .B1(new_n835_), .B2(new_n828_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n833_), .A2(new_n834_), .B1(new_n836_), .B2(KEYINPUT59), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n383_), .A2(G113gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n831_), .B1(new_n837_), .B2(new_n838_), .ZN(G1340gat));
  OAI21_X1  g638(.A(new_n834_), .B1(new_n832_), .B2(new_n828_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n830_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT121), .B1(new_n842_), .B2(new_n358_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n844_));
  INV_X1    g643(.A(new_n358_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n837_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n846_), .A3(G120gat), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n740_), .B2(G120gat), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n830_), .B(new_n849_), .C1(new_n848_), .C2(G120gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n830_), .B2(new_n231_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n852_), .A2(KEYINPUT122), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(KEYINPUT122), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n837_), .A2(G127gat), .A3(new_n627_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(G1342gat));
  AOI21_X1  g655(.A(G134gat), .B1(new_n830_), .B2(new_n736_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n813_), .A2(G134gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n837_), .B2(new_n858_), .ZN(G1343gat));
  NAND2_X1  g658(.A1(new_n825_), .A2(new_n829_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n513_), .ZN(new_n861_));
  AND4_X1   g660(.A1(new_n609_), .A2(new_n860_), .A3(new_n861_), .A4(new_n748_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n383_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n845_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT123), .B(G148gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1345gat));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n231_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT61), .B(G155gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT124), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n868_), .B(new_n870_), .ZN(G1346gat));
  AOI21_X1  g670(.A(G162gat), .B1(new_n862_), .B2(new_n736_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n813_), .A2(G162gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n862_), .B2(new_n873_), .ZN(G1347gat));
  NOR3_X1   g673(.A1(new_n748_), .A2(new_n609_), .A3(new_n515_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n833_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n376_), .B1(new_n876_), .B2(new_n383_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n833_), .A2(new_n875_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n878_), .A2(new_n551_), .A3(new_n826_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT62), .B1(new_n877_), .B2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G169gat), .B1(new_n878_), .B2(new_n826_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(G1348gat));
  AND2_X1   g683(.A1(new_n860_), .A2(new_n875_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(G176gat), .A3(new_n845_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n485_), .B1(new_n878_), .B2(new_n740_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n885_), .A2(KEYINPUT125), .A3(G176gat), .A4(new_n845_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(G1349gat));
  AOI21_X1  g690(.A(new_n473_), .B1(new_n885_), .B2(new_n231_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n229_), .A2(new_n553_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n876_), .B2(new_n893_), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n876_), .A2(new_n736_), .A3(new_n481_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G190gat), .B1(new_n878_), .B2(new_n684_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n896_), .A2(KEYINPUT126), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(KEYINPUT126), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n895_), .B1(new_n897_), .B2(new_n898_), .ZN(G1351gat));
  NOR2_X1   g698(.A1(new_n748_), .A2(new_n609_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n860_), .A2(new_n861_), .A3(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n378_), .B1(new_n901_), .B2(new_n826_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT127), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n901_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(G197gat), .A3(new_n383_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT127), .B(new_n378_), .C1(new_n901_), .C2(new_n826_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n904_), .A2(new_n906_), .A3(new_n907_), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n845_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n901_), .A2(new_n229_), .A3(new_n911_), .A4(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n905_), .A2(new_n627_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n911_), .ZN(G1354gat));
  INV_X1    g714(.A(G218gat), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n901_), .A2(new_n916_), .A3(new_n684_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n905_), .A2(new_n736_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n916_), .B2(new_n918_), .ZN(G1355gat));
endmodule


