//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n202_), .B(G43gat), .ZN(new_n206_));
  INV_X1    g005(.A(G50gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT79), .A2(G8gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT79), .A2(G8gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(G1gat), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT14), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n214_), .B2(KEYINPUT14), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n211_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G1gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(KEYINPUT14), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT80), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n216_), .ZN(new_n223_));
  INV_X1    g022(.A(G1gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n211_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n220_), .A2(new_n225_), .A3(G8gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(G8gat), .B1(new_n220_), .B2(new_n225_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n210_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n209_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n205_), .A2(new_n208_), .A3(KEYINPUT15), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G8gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n219_), .A2(G1gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n224_), .B1(new_n223_), .B2(new_n211_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n220_), .A2(new_n225_), .A3(G8gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n228_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT83), .B(G141gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(G169gat), .B(G197gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT82), .B(G113gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  NAND3_X1  g044(.A1(new_n236_), .A2(new_n209_), .A3(new_n237_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n228_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n240_), .B(new_n245_), .C1(new_n247_), .C2(new_n239_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n245_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n228_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n239_), .B1(new_n228_), .B2(new_n246_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n248_), .A2(new_n252_), .A3(KEYINPUT84), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT84), .B1(new_n248_), .B2(new_n252_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G99gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT10), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT10), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G99gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(new_n260_), .A3(KEYINPUT64), .ZN(new_n264_));
  AOI21_X1  g063(.A(G106gat), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n266_), .A2(KEYINPUT9), .ZN(new_n267_));
  NOR2_X1   g066(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(G92gat), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G85gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(G92gat), .ZN(new_n271_));
  INV_X1    g070(.A(G92gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(G85gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT9), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G99gat), .A2(G106gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT6), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(G99gat), .A3(G106gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n269_), .A2(new_n274_), .A3(new_n279_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n265_), .A2(new_n280_), .A3(KEYINPUT66), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282_));
  INV_X1    g081(.A(new_n279_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT9), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(KEYINPUT65), .A3(G85gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n270_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n272_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n272_), .A2(G85gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n270_), .A2(G92gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n284_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n283_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G106gat), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n258_), .A2(new_n260_), .A3(KEYINPUT64), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT64), .B1(new_n258_), .B2(new_n260_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n282_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT69), .B1(new_n281_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n257_), .A2(new_n293_), .A3(KEYINPUT67), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT7), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n301_), .A2(new_n257_), .A3(new_n293_), .A4(KEYINPUT67), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n279_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT8), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n289_), .A2(new_n290_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n276_), .A2(new_n278_), .A3(KEYINPUT68), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT68), .B1(new_n276_), .B2(new_n278_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n300_), .A2(new_n302_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n309_), .A2(new_n310_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n306_), .B1(new_n311_), .B2(new_n304_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT66), .B1(new_n265_), .B2(new_n280_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n288_), .A2(new_n291_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n296_), .A2(new_n282_), .A3(new_n314_), .A4(new_n279_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n298_), .A2(new_n312_), .A3(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G57gat), .B(G64gat), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(KEYINPUT11), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(KEYINPUT11), .ZN(new_n321_));
  XOR2_X1   g120(.A(G71gat), .B(G78gat), .Z(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n321_), .A2(new_n322_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT12), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n325_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n277_), .B1(G99gat), .B2(G106gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n275_), .A2(KEYINPUT6), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n276_), .A2(new_n278_), .A3(KEYINPUT68), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(new_n300_), .A3(new_n302_), .A4(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n305_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n329_), .B1(new_n336_), .B2(KEYINPUT8), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n313_), .A2(new_n315_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n328_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n318_), .A2(new_n327_), .B1(new_n339_), .B2(new_n326_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT70), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G230gat), .A2(G233gat), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n304_), .B1(new_n335_), .B2(new_n305_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n315_), .B(new_n313_), .C1(new_n343_), .C2(new_n329_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n341_), .B(new_n342_), .C1(new_n344_), .C2(new_n328_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n312_), .A2(new_n315_), .A3(new_n313_), .A4(new_n325_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n341_), .B1(new_n347_), .B2(new_n342_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n340_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n339_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(G230gat), .A3(G233gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G120gat), .B(G148gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G176gat), .B(G204gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n357_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n358_), .A2(KEYINPUT72), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT72), .B1(new_n358_), .B2(new_n359_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n363_));
  NAND2_X1  g162(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n364_));
  OR2_X1    g163(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n364_), .B(new_n365_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G127gat), .B(G134gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT88), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n368_), .B(new_n369_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n370_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT31), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(G183gat), .B2(G190gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n381_));
  OAI21_X1  g180(.A(G169gat), .B1(new_n381_), .B2(G176gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(G176gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(KEYINPUT85), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G169gat), .B(G176gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT25), .B(G183gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n387_), .A2(KEYINPUT24), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  OR3_X1    g189(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n379_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT86), .ZN(new_n394_));
  XOR2_X1   g193(.A(G71gat), .B(G99gat), .Z(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n394_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n398_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n374_), .B1(new_n403_), .B2(KEYINPUT89), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT87), .B1(new_n374_), .B2(KEYINPUT89), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT95), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT2), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT94), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n412_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(KEYINPUT92), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT3), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  NOR4_X1   g216(.A1(new_n417_), .A2(KEYINPUT92), .A3(G141gat), .A4(G148gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n414_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT93), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n408_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n415_), .B(KEYINPUT3), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n420_), .B(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n423_), .A2(KEYINPUT95), .A3(new_n414_), .A4(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n422_), .A2(new_n426_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n430_));
  OR3_X1    g229(.A1(new_n428_), .A2(new_n430_), .A3(KEYINPUT1), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(KEYINPUT1), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n428_), .B2(KEYINPUT1), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n431_), .A2(new_n427_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G141gat), .A2(G148gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n435_), .B(KEYINPUT90), .Z(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n436_), .A3(new_n409_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n429_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(KEYINPUT29), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G78gat), .B(G106gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G197gat), .A2(G204gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT96), .B(G197gat), .ZN(new_n444_));
  OAI211_X1 g243(.A(KEYINPUT21), .B(new_n443_), .C1(new_n444_), .C2(G204gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(G211gat), .B(G218gat), .Z(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G204gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G197gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n445_), .B(new_n447_), .C1(new_n450_), .C2(KEYINPUT21), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(KEYINPUT21), .A3(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n429_), .A2(new_n437_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT29), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n442_), .B(new_n453_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n429_), .B2(new_n437_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n453_), .ZN(new_n458_));
  OAI211_X1 g257(.A(G228gat), .B(G233gat), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G22gat), .B(G50gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT28), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n456_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n441_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n456_), .A2(new_n459_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n461_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n456_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n439_), .B(new_n440_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n438_), .A2(new_n373_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT101), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n454_), .A2(new_n372_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT101), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n438_), .A2(new_n477_), .A3(new_n373_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n475_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n479_), .A2(KEYINPUT4), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT4), .B1(new_n438_), .B2(new_n373_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n473_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n438_), .A2(new_n477_), .A3(new_n373_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n477_), .B1(new_n438_), .B2(new_n373_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT102), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n472_), .A4(new_n476_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n475_), .A2(new_n476_), .A3(new_n472_), .A4(new_n478_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT102), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT0), .B(G57gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G85gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(G1gat), .B(G29gat), .Z(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n482_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n481_), .B1(new_n479_), .B2(KEYINPUT4), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n487_), .B(new_n489_), .C1(new_n497_), .C2(new_n472_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n494_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n393_), .A2(new_n453_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT97), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT19), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT98), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n379_), .A2(new_n505_), .A3(new_n391_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n391_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT98), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n390_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G169gat), .A2(G176gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n383_), .A2(new_n384_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n380_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n509_), .A2(new_n512_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n513_));
  AND4_X1   g312(.A1(KEYINPUT20), .A2(new_n501_), .A3(new_n504_), .A4(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n512_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n453_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n392_), .A2(new_n386_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n504_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT18), .B(G64gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G92gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G8gat), .B(G36gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n524_), .A2(KEYINPUT32), .ZN(new_n525_));
  OR3_X1    g324(.A1(new_n514_), .A2(new_n519_), .A3(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n513_), .A2(KEYINPUT20), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n504_), .B1(new_n527_), .B2(new_n501_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n517_), .A2(new_n504_), .A3(new_n518_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n525_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n500_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT33), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n498_), .B2(new_n494_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n482_), .A2(new_n490_), .A3(KEYINPUT33), .A4(new_n495_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n519_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n527_), .A2(new_n504_), .A3(new_n501_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n524_), .A3(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n523_), .B1(new_n514_), .B2(new_n519_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(KEYINPUT99), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT100), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT99), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n535_), .A2(new_n541_), .A3(new_n536_), .A4(new_n524_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n539_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n485_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n494_), .B(new_n546_), .C1(new_n497_), .C2(new_n473_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n533_), .A2(new_n534_), .A3(new_n545_), .A4(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n471_), .B1(new_n531_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT27), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n539_), .A2(new_n550_), .A3(new_n542_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n523_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n537_), .A3(KEYINPUT27), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n471_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT103), .B1(new_n500_), .B2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n465_), .A2(new_n470_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n553_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT103), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(new_n499_), .A4(new_n496_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n407_), .B1(new_n549_), .B2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n407_), .A2(new_n500_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n557_), .A2(new_n471_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI211_X1 g364(.A(new_n256_), .B(new_n367_), .C1(new_n562_), .C2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT74), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT75), .B(KEYINPUT35), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n318_), .A2(new_n232_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT76), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n569_), .A2(new_n571_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n344_), .B2(new_n209_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n318_), .A2(KEYINPUT76), .A3(new_n232_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n576_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n572_), .A2(KEYINPUT78), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n579_), .A2(new_n574_), .A3(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n573_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n579_), .A2(new_n574_), .A3(new_n582_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(KEYINPUT78), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(KEYINPUT77), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(G134gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(G162gat), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n584_), .A2(KEYINPUT77), .A3(new_n587_), .A4(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n318_), .A2(KEYINPUT76), .A3(new_n232_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT76), .B1(new_n318_), .B2(new_n232_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n578_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n572_), .B1(new_n598_), .B2(new_n585_), .ZN(new_n599_));
  OAI211_X1 g398(.A(KEYINPUT36), .B(new_n591_), .C1(new_n599_), .C2(new_n586_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT16), .B(G183gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G211gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT81), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n226_), .A2(new_n227_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(new_n325_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n603_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n566_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n224_), .A3(new_n500_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT38), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n601_), .A2(KEYINPUT104), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n593_), .A2(new_n600_), .A3(new_n624_), .A4(new_n595_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n616_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n566_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n500_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n622_), .A2(new_n632_), .ZN(G1324gat));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n557_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G8gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT39), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n212_), .A2(new_n213_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n620_), .A2(new_n637_), .A3(new_n557_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g439(.A(G15gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n407_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n629_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT41), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n620_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n620_), .A2(new_n647_), .A3(new_n471_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G22gat), .B1(new_n630_), .B2(new_n556_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT105), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(KEYINPUT105), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(KEYINPUT42), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT42), .B1(new_n650_), .B2(new_n651_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n652_), .B2(new_n653_), .ZN(G1327gat));
  AOI21_X1  g453(.A(new_n626_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n367_), .A2(new_n617_), .A3(new_n256_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(G29gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n500_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n562_), .A2(new_n565_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n603_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT43), .B(new_n603_), .C1(new_n562_), .C2(new_n565_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n656_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT44), .B(new_n656_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(new_n500_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n659_), .B1(new_n670_), .B2(new_n658_), .ZN(G1328gat));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(KEYINPUT109), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n667_), .A2(new_n557_), .A3(new_n668_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT106), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n667_), .A2(new_n677_), .A3(new_n557_), .A4(new_n668_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(G36gat), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n676_), .A2(KEYINPUT107), .A3(G36gat), .A4(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n672_), .A2(KEYINPUT109), .ZN(new_n684_));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n657_), .A2(new_n685_), .A3(new_n557_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT108), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n657_), .A2(new_n689_), .A3(new_n685_), .A4(new_n557_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n687_), .A2(new_n688_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n688_), .B1(new_n687_), .B2(new_n690_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n684_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n674_), .B1(new_n683_), .B2(new_n694_), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n673_), .B(new_n693_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  NAND3_X1  g496(.A1(new_n669_), .A2(G43gat), .A3(new_n642_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n657_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n203_), .B1(new_n699_), .B2(new_n407_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g501(.A1(new_n657_), .A2(new_n207_), .A3(new_n471_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n669_), .A2(new_n471_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n704_), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT110), .B1(new_n704_), .B2(G50gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(G1331gat));
  AND3_X1   g506(.A1(new_n661_), .A2(new_n256_), .A3(new_n367_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n628_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(G57gat), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n631_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n619_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(KEYINPUT111), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(KEYINPUT111), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n500_), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n716_), .B2(new_n711_), .ZN(G1332gat));
  INV_X1    g516(.A(G64gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n709_), .B2(new_n557_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT48), .Z(new_n720_));
  INV_X1    g519(.A(new_n713_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n718_), .A3(new_n557_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1333gat));
  OR3_X1    g522(.A1(new_n713_), .A2(G71gat), .A3(new_n407_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G71gat), .B1(new_n710_), .B2(new_n407_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT112), .Z(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT49), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT49), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n709_), .B2(new_n471_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT50), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n721_), .A2(new_n730_), .A3(new_n471_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1335gat));
  INV_X1    g533(.A(new_n367_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n735_), .A2(new_n617_), .A3(new_n255_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n655_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n270_), .B1(new_n737_), .B2(new_n631_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n663_), .A2(new_n664_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n736_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT113), .Z(new_n741_));
  INV_X1    g540(.A(new_n266_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n500_), .B1(new_n268_), .B2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n738_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT114), .Z(G1336gat));
  INV_X1    g544(.A(new_n737_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G92gat), .B1(new_n746_), .B2(new_n557_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n741_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n272_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(G1337gat));
  OAI21_X1  g549(.A(G99gat), .B1(new_n741_), .B2(new_n407_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n407_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT115), .B1(new_n746_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g554(.A(G106gat), .B1(new_n740_), .B2(new_n556_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT52), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n746_), .A2(new_n293_), .A3(new_n471_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g559(.A(G113gat), .ZN(new_n761_));
  INV_X1    g560(.A(new_n239_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n228_), .A2(new_n238_), .A3(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n249_), .B(new_n763_), .C1(new_n247_), .C2(new_n762_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(new_n248_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n340_), .B(KEYINPUT55), .C1(new_n348_), .C2(new_n346_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n340_), .A2(new_n347_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(G230gat), .A3(G233gat), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n772_));
  NAND2_X1  g571(.A1(new_n349_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n342_), .B1(new_n344_), .B2(new_n328_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT70), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n345_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n340_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n769_), .A2(new_n771_), .A3(new_n773_), .A4(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n357_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n358_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT118), .B1(new_n778_), .B2(new_n357_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n255_), .B1(new_n783_), .B2(KEYINPUT56), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n766_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(KEYINPUT57), .A3(new_n626_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT121), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n785_), .A2(new_n626_), .A3(new_n788_), .A4(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n785_), .A2(new_n626_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n357_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT119), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n778_), .A2(new_n797_), .A3(KEYINPUT56), .A4(new_n357_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n778_), .C2(new_n357_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n779_), .B2(new_n802_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n799_), .A2(new_n800_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n765_), .A2(new_n358_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n794_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n805_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n803_), .A2(new_n800_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT58), .B(new_n807_), .C1(new_n808_), .C2(new_n799_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n809_), .A3(new_n662_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n790_), .A2(new_n793_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT122), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n790_), .A2(new_n793_), .A3(new_n810_), .A4(KEYINPUT122), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n616_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n618_), .A2(new_n367_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n256_), .ZN(new_n818_));
  NOR4_X1   g617(.A1(new_n618_), .A2(new_n367_), .A3(KEYINPUT54), .A4(new_n255_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n815_), .A2(new_n821_), .ZN(new_n822_));
  NOR4_X1   g621(.A1(new_n407_), .A2(new_n631_), .A3(new_n471_), .A4(new_n557_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n761_), .B1(new_n824_), .B2(new_n256_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n811_), .A2(new_n828_), .A3(new_n616_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n811_), .B2(new_n616_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n820_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n823_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n827_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n811_), .A2(new_n616_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT123), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n811_), .A2(new_n828_), .A3(new_n616_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n821_), .A3(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(KEYINPUT124), .A3(new_n832_), .A4(new_n823_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n826_), .A2(new_n834_), .A3(G113gat), .A4(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n825_), .B1(new_n840_), .B2(new_n256_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT125), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n825_), .B(new_n843_), .C1(new_n840_), .C2(new_n256_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1340gat));
  INV_X1    g644(.A(new_n824_), .ZN(new_n846_));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n735_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n846_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  AND4_X1   g648(.A1(new_n367_), .A2(new_n826_), .A3(new_n834_), .A4(new_n839_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n847_), .ZN(G1341gat));
  AOI21_X1  g650(.A(G127gat), .B1(new_n846_), .B2(new_n617_), .ZN(new_n852_));
  AND4_X1   g651(.A1(new_n617_), .A2(new_n826_), .A3(new_n834_), .A4(new_n839_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g653(.A(G134gat), .B1(new_n846_), .B2(new_n627_), .ZN(new_n855_));
  AND4_X1   g654(.A1(new_n662_), .A2(new_n826_), .A3(new_n834_), .A4(new_n839_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(G134gat), .ZN(G1343gat));
  AOI21_X1  g656(.A(new_n642_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n858_), .A2(new_n500_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(new_n255_), .A3(new_n558_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n558_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n735_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT126), .B(G148gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1345gat));
  NOR2_X1   g664(.A1(new_n862_), .A2(new_n616_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT61), .B(G155gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  INV_X1    g667(.A(G162gat), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n862_), .A2(new_n869_), .A3(new_n603_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n859_), .A2(new_n627_), .A3(new_n558_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(new_n871_), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n831_), .A2(new_n471_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n563_), .A2(new_n557_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n255_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G169gat), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n873_), .A2(new_n874_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n255_), .A3(new_n383_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n875_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(G1348gat));
  AOI21_X1  g681(.A(G176gat), .B1(new_n879_), .B2(new_n367_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n471_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n884_), .A2(G176gat), .A3(new_n367_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n874_), .B2(new_n885_), .ZN(G1349gat));
  NAND2_X1  g685(.A1(new_n874_), .A2(new_n617_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G183gat), .B1(new_n884_), .B2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n388_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n873_), .B2(new_n890_), .ZN(G1350gat));
  NAND2_X1  g690(.A1(new_n879_), .A2(new_n662_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G190gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n879_), .A2(new_n627_), .A3(new_n389_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1351gat));
  AOI21_X1  g694(.A(new_n500_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n858_), .A2(new_n471_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n255_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n367_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n903_));
  INV_X1    g702(.A(G211gat), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n897_), .A2(new_n902_), .A3(new_n617_), .A4(new_n906_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n858_), .A2(new_n617_), .A3(new_n471_), .A4(new_n896_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT127), .B1(new_n908_), .B2(new_n905_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n903_), .A2(new_n904_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n907_), .A2(new_n903_), .A3(new_n909_), .A4(new_n904_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1354gat));
  AOI21_X1  g713(.A(G218gat), .B1(new_n897_), .B2(new_n627_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n897_), .A2(new_n662_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(G218gat), .B2(new_n916_), .ZN(G1355gat));
endmodule


