//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT88), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n204_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n211_), .A2(new_n204_), .A3(new_n214_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n207_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(new_n210_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT22), .B(G169gat), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT89), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT89), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(G176gat), .B1(new_n225_), .B2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n220_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n208_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT90), .B1(new_n229_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n228_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n226_), .A2(new_n227_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n206_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT90), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n220_), .A2(new_n230_), .B1(G169gat), .B2(G176gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n218_), .A2(new_n223_), .B1(new_n233_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G211gat), .B(G218gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT21), .ZN(new_n244_));
  OR2_X1    g043(.A1(G197gat), .A2(G204gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G197gat), .A2(G204gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n243_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT85), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n241_), .A2(new_n242_), .ZN(new_n250_));
  INV_X1    g049(.A(G218gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G211gat), .ZN(new_n252_));
  INV_X1    g051(.A(G211gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G218gat), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n252_), .A2(new_n254_), .A3(new_n242_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT83), .B1(new_n245_), .B2(new_n246_), .ZN(new_n256_));
  OAI22_X1  g055(.A1(new_n250_), .A2(new_n255_), .B1(new_n244_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n244_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n249_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n256_), .A2(new_n244_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n243_), .A2(new_n261_), .A3(KEYINPUT85), .A4(new_n258_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n248_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT20), .B1(new_n240_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n262_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n248_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G183gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT73), .B1(new_n268_), .B2(KEYINPUT25), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n269_), .B(new_n213_), .C1(new_n212_), .C2(KEYINPUT73), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n209_), .B2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n207_), .A2(KEYINPUT74), .A3(KEYINPUT24), .A4(new_n208_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT75), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n270_), .A2(new_n273_), .A3(new_n277_), .A4(new_n274_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n221_), .B1(new_n272_), .B2(new_n222_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n281_));
  NAND2_X1  g080(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n205_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT77), .ZN(new_n284_));
  AOI21_X1  g083(.A(G176gat), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT77), .B1(new_n205_), .B2(KEYINPUT22), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT78), .B1(new_n220_), .B2(new_n230_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n220_), .A2(KEYINPUT78), .A3(new_n230_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n287_), .B(new_n208_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n280_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n267_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n203_), .B1(new_n264_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n267_), .A2(new_n291_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT20), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n203_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n233_), .A2(new_n239_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n211_), .A2(new_n204_), .A3(new_n214_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n223_), .B1(new_n298_), .B2(new_n215_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n294_), .B(new_n296_), .C1(new_n267_), .C2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT18), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT91), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n293_), .A2(new_n301_), .A3(new_n307_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT27), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT97), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n299_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT20), .B1(new_n315_), .B2(new_n267_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n263_), .B1(new_n290_), .B2(new_n280_), .ZN(new_n317_));
  OAI211_X1 g116(.A(KEYINPUT96), .B(new_n203_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n295_), .B1(new_n300_), .B2(new_n267_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n203_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n319_), .B(new_n320_), .C1(new_n291_), .C2(new_n267_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n294_), .B(KEYINPUT20), .C1(new_n267_), .C2(new_n315_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT96), .B1(new_n323_), .B2(new_n203_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n308_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n293_), .A2(KEYINPUT97), .A3(new_n301_), .A4(new_n307_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n314_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT98), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT98), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n314_), .A2(new_n325_), .A3(new_n329_), .A4(new_n326_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n311_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  OR2_X1    g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n335_), .B(KEYINPUT3), .Z(new_n336_));
  NAND2_X1  g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT2), .Z(new_n338_));
  OAI211_X1 g137(.A(new_n333_), .B(new_n334_), .C1(new_n336_), .C2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n335_), .B(KEYINPUT80), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n342_), .A2(new_n333_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n333_), .A2(KEYINPUT1), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n337_), .B(new_n340_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G113gat), .B(G120gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT92), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT92), .ZN(new_n353_));
  INV_X1    g152(.A(new_n347_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n354_), .A2(new_n348_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n348_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT79), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n349_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n353_), .B1(new_n360_), .B2(new_n346_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n352_), .B(KEYINPUT4), .C1(new_n351_), .C2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n346_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT4), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n332_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n346_), .A2(new_n353_), .A3(new_n350_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(KEYINPUT92), .ZN(new_n367_));
  INV_X1    g166(.A(new_n351_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n332_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G57gat), .B(G85gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT94), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT93), .B(KEYINPUT0), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  OR3_X1    g176(.A1(new_n365_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n365_), .B2(new_n371_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n280_), .A2(new_n290_), .A3(KEYINPUT30), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383_));
  INV_X1    g182(.A(G43gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(G15gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n385_), .B(new_n388_), .Z(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT30), .B1(new_n280_), .B2(new_n290_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n382_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n291_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n389_), .B1(new_n394_), .B2(new_n381_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT31), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n390_), .B1(new_n382_), .B2(new_n391_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT31), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n389_), .A3(new_n381_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n360_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n360_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n339_), .A2(new_n345_), .A3(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G22gat), .B(G50gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n404_), .B1(new_n339_), .B2(new_n345_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n267_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n408_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n263_), .B2(new_n409_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT86), .Z(new_n415_));
  AND3_X1   g214(.A1(new_n411_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n407_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(KEYINPUT28), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT82), .ZN(new_n420_));
  INV_X1    g219(.A(new_n415_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n408_), .B1(new_n267_), .B2(new_n410_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n263_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n407_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n411_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n418_), .A2(new_n420_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n420_), .B1(new_n418_), .B2(new_n427_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n401_), .B(new_n403_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n420_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n416_), .A2(new_n417_), .A3(new_n407_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n425_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n418_), .A2(new_n420_), .A3(new_n427_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n401_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n434_), .B(new_n435_), .C1(new_n436_), .C2(new_n402_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n380_), .B1(new_n430_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n307_), .A2(KEYINPUT32), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n322_), .A2(new_n324_), .A3(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n302_), .A2(new_n439_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n380_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(KEYINPUT33), .B(new_n377_), .C1(new_n365_), .C2(new_n371_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT95), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n379_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n377_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n370_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n369_), .A2(new_n332_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n447_), .A2(new_n310_), .A3(new_n309_), .A4(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n442_), .B1(new_n445_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n428_), .A2(new_n429_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n436_), .A2(new_n402_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n331_), .A2(new_n438_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G99gat), .ZN(new_n461_));
  INV_X1    g260(.A(G106gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT64), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT7), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT7), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(new_n461_), .A3(new_n462_), .A4(KEYINPUT64), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n460_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G85gat), .B(G92gat), .Z(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT65), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(KEYINPUT65), .A3(new_n468_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT8), .A3(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G57gat), .B(G64gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G71gat), .B(G78gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n476_), .B1(KEYINPUT11), .B2(new_n474_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT8), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n469_), .A2(new_n470_), .A3(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT10), .B(G99gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n462_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n468_), .A2(KEYINPUT9), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT9), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(G85gat), .A3(G92gat), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n486_), .A2(new_n487_), .A3(new_n460_), .A4(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n473_), .A2(new_n482_), .A3(new_n484_), .A4(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G230gat), .A2(G233gat), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT12), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n472_), .A2(KEYINPUT8), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT65), .B1(new_n467_), .B2(new_n468_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n490_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n484_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n494_), .B(new_n481_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n473_), .A2(new_n484_), .A3(new_n490_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n494_), .B1(new_n501_), .B2(new_n481_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n493_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT66), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n481_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n491_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n492_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT66), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n509_), .B(new_n493_), .C1(new_n500_), .C2(new_n502_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n504_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G120gat), .B(G148gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT5), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G176gat), .B(G204gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n504_), .A2(new_n508_), .A3(new_n510_), .A4(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT13), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521_));
  INV_X1    g320(.A(G1gat), .ZN(new_n522_));
  INV_X1    g321(.A(G8gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G1gat), .B(G8gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G29gat), .B(G36gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(new_n531_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(KEYINPUT70), .A3(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(KEYINPUT70), .B2(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n530_), .B(KEYINPUT15), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n532_), .B1(new_n539_), .B2(new_n527_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n537_), .B(KEYINPUT71), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G113gat), .B(G141gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT72), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n538_), .A2(new_n542_), .A3(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n520_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n501_), .A2(new_n539_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT68), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n473_), .A2(new_n530_), .A3(new_n484_), .A4(new_n490_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G190gat), .B(G218gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n560_), .A2(new_n563_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n564_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n567_), .B(KEYINPUT36), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(KEYINPUT69), .A2(KEYINPUT37), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n572_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT69), .B(KEYINPUT37), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n564_), .A2(new_n570_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n573_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n581_), .B2(new_n571_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n527_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n481_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT16), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n587_), .A2(new_n588_), .A3(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(KEYINPUT17), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n583_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n457_), .A2(new_n552_), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT99), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n522_), .A3(new_n380_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n331_), .A2(new_n438_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n453_), .A2(new_n456_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n581_), .A2(KEYINPUT102), .A3(new_n571_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(new_n597_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n552_), .A2(KEYINPUT101), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n519_), .A2(KEYINPUT13), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT13), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n613_), .B(new_n551_), .C1(new_n614_), .C2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n611_), .B1(new_n612_), .B2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(new_n380_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n603_), .B1(new_n522_), .B2(new_n619_), .ZN(G1324gat));
  INV_X1    g419(.A(new_n331_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n600_), .A2(new_n523_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT103), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n523_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT39), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1325gat));
  INV_X1    g427(.A(new_n455_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n387_), .B1(new_n618_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n600_), .A2(new_n387_), .A3(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n454_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n618_), .B2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n600_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n610_), .A2(new_n597_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n457_), .A2(new_n552_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n380_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n597_), .B1(new_n612_), .B2(new_n617_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  INV_X1    g445(.A(new_n583_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n606_), .B2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n457_), .A2(KEYINPUT43), .A3(new_n583_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT44), .B(new_n645_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n650_), .A2(G29gat), .A3(new_n380_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n648_), .A2(new_n649_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n613_), .B1(new_n520_), .B2(new_n551_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n617_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n596_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n644_), .B1(new_n651_), .B2(new_n657_), .ZN(G1328gat));
  INV_X1    g457(.A(new_n552_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n606_), .A2(new_n659_), .A3(new_n641_), .ZN(new_n660_));
  INV_X1    g459(.A(G36gat), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n331_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n331_), .A2(new_n662_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT108), .B1(new_n660_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n621_), .A2(KEYINPUT106), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n331_), .A2(new_n662_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G36gat), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT108), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n643_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n666_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n666_), .B2(new_n671_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n650_), .A2(new_n621_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n606_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n457_), .B2(new_n583_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n656_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(KEYINPUT44), .ZN(new_n681_));
  OAI21_X1  g480(.A(G36gat), .B1(new_n677_), .B2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT110), .B1(new_n676_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT111), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT110), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n331_), .B1(new_n680_), .B2(KEYINPUT44), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n661_), .B1(new_n687_), .B2(new_n657_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n666_), .A2(new_n671_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n672_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n666_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n686_), .B1(new_n688_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(KEYINPUT46), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT109), .B1(new_n676_), .B2(new_n682_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n686_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n685_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n685_), .B2(new_n695_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  OAI21_X1  g499(.A(new_n384_), .B1(new_n660_), .B2(new_n455_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n650_), .A2(G43gat), .A3(new_n629_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n681_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(G1330gat));
  AOI21_X1  g504(.A(G50gat), .B1(new_n643_), .B2(new_n635_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n650_), .A2(G50gat), .A3(new_n635_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n657_), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n520_), .A2(new_n551_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n710_), .A2(new_n457_), .A3(new_n598_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n380_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n606_), .A2(new_n597_), .A3(new_n610_), .A4(new_n709_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT113), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n380_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n716_), .B2(new_n712_), .ZN(G1332gat));
  INV_X1    g516(.A(G64gat), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n667_), .A2(new_n668_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n715_), .B2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT48), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n711_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1333gat));
  INV_X1    g522(.A(G71gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n715_), .B2(new_n629_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT49), .Z(new_n726_));
  NAND3_X1  g525(.A1(new_n711_), .A2(new_n724_), .A3(new_n629_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1334gat));
  INV_X1    g527(.A(G78gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n715_), .B2(new_n635_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT50), .Z(new_n731_));
  NAND3_X1  g530(.A1(new_n711_), .A2(new_n729_), .A3(new_n635_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1335gat));
  OAI211_X1 g532(.A(new_n596_), .B(new_n709_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT115), .ZN(new_n735_));
  INV_X1    g534(.A(G85gat), .ZN(new_n736_));
  INV_X1    g535(.A(new_n380_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n710_), .A2(new_n457_), .A3(new_n642_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n380_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT114), .Z(new_n741_));
  NOR2_X1   g540(.A1(new_n738_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT116), .ZN(G1336gat));
  NAND2_X1  g542(.A1(new_n719_), .A2(G92gat), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT117), .Z(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n739_), .A2(new_n621_), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n735_), .A2(new_n746_), .B1(G92gat), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT118), .ZN(G1337gat));
  NAND3_X1  g548(.A1(new_n739_), .A2(new_n485_), .A3(new_n629_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n735_), .A2(new_n455_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n461_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n739_), .A2(new_n462_), .A3(new_n635_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G106gat), .B1(new_n734_), .B2(new_n454_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT52), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT52), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g558(.A1(new_n551_), .A2(new_n596_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT119), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n614_), .A2(new_n616_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n647_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n763_), .A2(new_n764_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n551_), .A2(new_n518_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n504_), .A2(new_n771_), .A3(new_n510_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n491_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n491_), .A2(new_n492_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n505_), .A2(KEYINPUT12), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n499_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n507_), .A2(new_n773_), .B1(new_n776_), .B2(KEYINPUT55), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n772_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n515_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n515_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n770_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n541_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n547_), .B1(new_n540_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n536_), .B2(new_n784_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n550_), .A2(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n519_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n610_), .B1(new_n783_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n787_), .A2(new_n518_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n515_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n780_), .B(new_n517_), .C1(new_n772_), .C2(new_n777_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n583_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n781_), .A2(new_n782_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n792_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n792_), .B(KEYINPUT58), .C1(new_n793_), .C2(new_n794_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n797_), .A2(new_n799_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n791_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n789_), .A2(new_n790_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n596_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n769_), .A2(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n621_), .A2(new_n737_), .A3(new_n437_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810_), .B2(new_n551_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n804_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n805_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n791_), .A2(new_n803_), .A3(KEYINPUT121), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n816_), .A2(KEYINPUT122), .A3(new_n596_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT122), .B1(new_n816_), .B2(new_n596_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n769_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n808_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n819_), .A2(new_n822_), .B1(new_n809_), .B2(KEYINPUT59), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n551_), .A2(new_n824_), .A3(G113gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n824_), .B2(G113gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n811_), .B1(new_n823_), .B2(new_n826_), .ZN(G1340gat));
  NAND2_X1  g626(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n791_), .A2(new_n803_), .A3(KEYINPUT121), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT121), .B1(new_n791_), .B2(new_n803_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n805_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n832_), .B2(new_n597_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n816_), .A2(KEYINPUT122), .A3(new_n596_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n768_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n762_), .B(new_n828_), .C1(new_n835_), .C2(new_n821_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT124), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n819_), .A2(new_n822_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n762_), .A4(new_n828_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(G120gat), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n842_));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n762_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n810_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n841_), .A2(new_n846_), .ZN(G1341gat));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n810_), .A2(new_n848_), .A3(new_n597_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n823_), .A2(new_n597_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n848_), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  INV_X1    g651(.A(new_n610_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n810_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n823_), .A2(new_n647_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n852_), .ZN(G1343gat));
  AOI21_X1  g655(.A(new_n430_), .B1(new_n769_), .B2(new_n806_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n719_), .A2(new_n737_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n551_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n762_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g663(.A1(new_n859_), .A2(new_n596_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT61), .B(G155gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  OR3_X1    g666(.A1(new_n859_), .A2(G162gat), .A3(new_n610_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G162gat), .B1(new_n859_), .B2(new_n583_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1347gat));
  AOI21_X1  g669(.A(new_n380_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n629_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT125), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n635_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n819_), .A2(new_n551_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G169gat), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n234_), .A2(new_n235_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n878_), .B(new_n879_), .C1(new_n880_), .C2(new_n875_), .ZN(G1348gat));
  NOR3_X1   g680(.A1(new_n835_), .A2(new_n635_), .A3(new_n873_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G176gat), .B1(new_n882_), .B2(new_n762_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n635_), .B1(new_n769_), .B2(new_n806_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n873_), .A2(new_n206_), .A3(new_n520_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1349gat));
  NOR2_X1   g685(.A1(new_n873_), .A2(new_n596_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G183gat), .B1(new_n887_), .B2(new_n884_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n596_), .A2(new_n212_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n882_), .B2(new_n889_), .ZN(G1350gat));
  NAND2_X1  g689(.A1(new_n882_), .A2(new_n647_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G190gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n882_), .A2(new_n213_), .A3(new_n853_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1351gat));
  NAND2_X1  g693(.A1(new_n857_), .A2(new_n871_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n551_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n762_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g699(.A(new_n596_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n901_), .B(KEYINPUT126), .Z(new_n902_));
  NAND2_X1  g701(.A1(new_n896_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n903_), .B(new_n904_), .Z(G1354gat));
  OAI21_X1  g704(.A(G218gat), .B1(new_n895_), .B2(new_n583_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n853_), .A2(new_n251_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n895_), .B2(new_n907_), .ZN(G1355gat));
endmodule


