//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(new_n204_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n208_), .A3(new_n206_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT88), .ZN(new_n213_));
  INV_X1    g012(.A(G155gat), .ZN(new_n214_));
  INV_X1    g013(.A(G162gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n214_), .A2(new_n215_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G141gat), .ZN(new_n221_));
  INV_X1    g020(.A(G148gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT90), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(new_n227_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n224_), .A2(KEYINPUT2), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G141gat), .A3(G148gat), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n234_), .A2(new_n236_), .B1(new_n223_), .B2(KEYINPUT3), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(new_n233_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT88), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n212_), .B(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(new_n217_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT91), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n238_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n226_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT29), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n211_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G228gat), .ZN(new_n249_));
  INV_X1    g048(.A(G233gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n238_), .A2(new_n244_), .A3(new_n241_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n244_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n225_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n210_), .B1(new_n255_), .B2(KEYINPUT29), .ZN(new_n256_));
  INV_X1    g055(.A(new_n251_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G78gat), .B(G106gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT92), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n252_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n202_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n246_), .A2(new_n266_), .A3(new_n247_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT28), .B1(new_n255_), .B2(KEYINPUT29), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G22gat), .B(G50gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n268_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n261_), .B1(new_n252_), .B2(new_n258_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n270_), .B(new_n273_), .C1(new_n274_), .C2(KEYINPUT93), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT94), .B1(new_n265_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n270_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n263_), .B2(new_n202_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n264_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT93), .B1(new_n279_), .B2(new_n274_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT94), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n277_), .B1(new_n279_), .B2(new_n274_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT22), .B(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n287_), .A2(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n292_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n291_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT82), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(G169gat), .B2(G176gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n299_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n288_), .A2(new_n287_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT25), .B(G183gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT26), .B(G190gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n303_), .A3(new_n299_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n292_), .A2(KEYINPUT85), .A3(new_n293_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT85), .B1(new_n295_), .B2(new_n292_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n292_), .A2(new_n293_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n298_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT86), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(new_n298_), .C1(new_n311_), .C2(new_n315_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n210_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n289_), .A2(new_n290_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n305_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT96), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n291_), .A2(KEYINPUT96), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n329_), .B(new_n330_), .C1(new_n315_), .C2(new_n297_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n296_), .B1(new_n304_), .B2(new_n286_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n300_), .A2(new_n299_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n309_), .A3(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n210_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n321_), .A2(KEYINPUT20), .A3(new_n325_), .A4(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT20), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n331_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n211_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n317_), .A2(new_n210_), .A3(new_n319_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n324_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344_));
  INV_X1    g143(.A(G92gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT18), .B(G64gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n337_), .A2(new_n343_), .A3(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n342_), .A2(new_n324_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n321_), .A2(KEYINPUT20), .A3(new_n336_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n324_), .B2(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n348_), .B(KEYINPUT100), .Z(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT27), .B(new_n350_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  NOR4_X1   g154(.A1(new_n320_), .A2(new_n335_), .A3(new_n338_), .A4(new_n324_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n325_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n348_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n350_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  INV_X1    g162(.A(G120gat), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n364_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT87), .B(G113gat), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G227gat), .A2(G233gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(KEYINPUT31), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n370_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n317_), .A2(new_n319_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G43gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT30), .B(G15gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n375_), .B(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n370_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n255_), .A2(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n370_), .B(new_n225_), .C1(new_n254_), .C2(new_n253_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(KEYINPUT4), .A3(new_n386_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n255_), .A2(new_n389_), .A3(new_n384_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n391_), .B2(new_n383_), .ZN(new_n392_));
  XOR2_X1   g191(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n393_));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n392_), .A2(new_n398_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n381_), .A2(new_n401_), .ZN(new_n402_));
  OR3_X1    g201(.A1(new_n285_), .A2(new_n362_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT98), .B1(new_n392_), .B2(new_n398_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT33), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n385_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n398_), .B(new_n406_), .C1(new_n391_), .C2(new_n383_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n358_), .A2(new_n407_), .A3(new_n350_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT98), .B(new_n409_), .C1(new_n392_), .C2(new_n398_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT99), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n337_), .A2(new_n343_), .A3(new_n413_), .ZN(new_n414_));
  OAI221_X1 g213(.A(new_n414_), .B1(new_n353_), .B2(new_n413_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n405_), .A2(new_n408_), .A3(new_n416_), .A4(new_n410_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n412_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n285_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n401_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n362_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n418_), .A2(new_n419_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n403_), .B1(new_n423_), .B2(new_n381_), .ZN(new_n424_));
  INV_X1    g223(.A(G1gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT75), .B(G8gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT14), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G15gat), .B(G22gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n425_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n428_), .A2(new_n430_), .A3(new_n425_), .ZN(new_n431_));
  OR3_X1    g230(.A1(new_n429_), .A2(new_n431_), .A3(G8gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(G8gat), .B1(new_n429_), .B2(new_n431_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(G231gat), .B2(G233gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G231gat), .A2(G233gat), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT68), .B(G71gat), .ZN(new_n439_));
  INV_X1    g238(.A(G78gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G57gat), .B(G64gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n439_), .A2(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n439_), .A2(new_n440_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n443_), .A4(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n438_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n457_));
  XNOR2_X1  g256(.A(G127gat), .B(G155gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G183gat), .B(G211gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n461_), .A2(KEYINPUT17), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(KEYINPUT17), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n452_), .A2(new_n453_), .A3(KEYINPUT78), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n456_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n454_), .A2(new_n462_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n454_), .A2(KEYINPUT77), .A3(new_n462_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  INV_X1    g272(.A(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT10), .B(G99gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n480_), .B2(new_n475_), .ZN(new_n481_));
  AND2_X1   g280(.A1(G85gat), .A2(G92gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G85gat), .A2(G92gat), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n482_), .A2(new_n483_), .B1(KEYINPUT64), .B2(KEYINPUT9), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n486_));
  NOR2_X1   g285(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n484_), .A2(new_n488_), .A3(KEYINPUT65), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT65), .B1(new_n484_), .B2(new_n488_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n481_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT66), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT66), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n481_), .B(new_n493_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n494_));
  OR3_X1    g293(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n495_), .A2(new_n476_), .A3(new_n477_), .A4(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n482_), .A2(new_n483_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT67), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT8), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n497_), .A2(new_n500_), .A3(new_n501_), .A4(new_n498_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n492_), .A2(new_n494_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT15), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT34), .ZN(new_n513_));
  INV_X1    g312(.A(new_n509_), .ZN(new_n514_));
  OAI221_X1 g313(.A(new_n511_), .B1(KEYINPUT35), .B2(new_n513_), .C1(new_n514_), .C2(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(KEYINPUT35), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  XNOR2_X1  g316(.A(G190gat), .B(G218gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(new_n215_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT73), .B(G134gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT36), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(KEYINPUT36), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n517_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n515_), .B(new_n516_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT74), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n530_), .A3(KEYINPUT37), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT37), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n525_), .B(new_n527_), .C1(new_n529_), .C2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n424_), .A2(new_n472_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT79), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n432_), .A2(new_n433_), .A3(new_n509_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n509_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n537_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(KEYINPUT79), .A3(new_n538_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n536_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n434_), .A2(new_n510_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n545_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT80), .B(G113gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G141gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G169gat), .B(G197gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  OR3_X1    g349(.A1(new_n544_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT81), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(KEYINPUT81), .B(new_n550_), .C1(new_n544_), .C2(new_n546_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n506_), .A2(new_n451_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n506_), .A2(new_n451_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT69), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n492_), .A2(new_n450_), .A3(new_n494_), .A4(new_n505_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n566_), .A2(KEYINPUT70), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT70), .B1(new_n566_), .B2(new_n567_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n560_), .B(new_n565_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n561_), .A2(new_n566_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G176gat), .B(G204gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n570_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n580_), .A2(KEYINPUT13), .A3(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT13), .B1(new_n580_), .B2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT72), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n535_), .A2(new_n557_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT101), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n425_), .A3(new_n420_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n584_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n556_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n424_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n472_), .A3(new_n528_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n401_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n589_), .A2(new_n590_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(new_n596_), .A3(new_n597_), .ZN(G1324gat));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n426_), .A3(new_n362_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G8gat), .B1(new_n595_), .B2(new_n422_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT39), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g402(.A(G15gat), .B1(new_n595_), .B2(new_n380_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT103), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT41), .ZN(new_n606_));
  INV_X1    g405(.A(G15gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n588_), .A2(new_n607_), .A3(new_n381_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(G1326gat));
  INV_X1    g408(.A(G22gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n588_), .A2(new_n610_), .A3(new_n285_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G22gat), .B1(new_n595_), .B2(new_n419_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT42), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(G1327gat));
  INV_X1    g413(.A(KEYINPUT105), .ZN(new_n615_));
  INV_X1    g414(.A(new_n534_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n418_), .A2(new_n419_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n421_), .A2(new_n422_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n381_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n403_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n615_), .B(new_n616_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT104), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT43), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT105), .B(new_n403_), .C1(new_n423_), .C2(new_n381_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n471_), .B1(new_n624_), .B2(new_n534_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n424_), .A2(new_n616_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT43), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(KEYINPUT104), .A3(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n623_), .A2(new_n593_), .A3(new_n626_), .A4(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT106), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n401_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(G29gat), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n472_), .A2(new_n528_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n594_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n420_), .A2(new_n636_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT107), .ZN(new_n640_));
  OAI22_X1  g439(.A1(new_n635_), .A2(new_n636_), .B1(new_n638_), .B2(new_n640_), .ZN(G1328gat));
  NOR3_X1   g440(.A1(new_n638_), .A2(G36gat), .A3(new_n422_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n422_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n645_));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT46), .B(new_n644_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1329gat));
  INV_X1    g450(.A(KEYINPUT47), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n630_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT44), .B1(new_n630_), .B2(KEYINPUT106), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n381_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G43gat), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n638_), .A2(G43gat), .A3(new_n380_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n652_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT47), .B(new_n657_), .C1(new_n655_), .C2(G43gat), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1330gat));
  INV_X1    g460(.A(G50gat), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n594_), .A2(new_n662_), .A3(new_n285_), .A4(new_n637_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n419_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(new_n662_), .ZN(G1331gat));
  NOR2_X1   g464(.A1(new_n557_), .A2(new_n471_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n424_), .A2(new_n528_), .A3(new_n585_), .A4(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT109), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(G57gat), .A3(new_n420_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT110), .Z(new_n670_));
  NOR2_X1   g469(.A1(new_n584_), .A2(new_n557_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n535_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G57gat), .B1(new_n672_), .B2(new_n420_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n670_), .A2(new_n673_), .ZN(G1332gat));
  INV_X1    g473(.A(G64gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n668_), .B2(new_n362_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT48), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n672_), .A2(new_n675_), .A3(new_n362_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1333gat));
  INV_X1    g478(.A(G71gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n668_), .B2(new_n381_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT49), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n672_), .A2(new_n680_), .A3(new_n381_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1334gat));
  NAND3_X1  g483(.A1(new_n672_), .A2(new_n440_), .A3(new_n285_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT50), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n668_), .A2(new_n285_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(G78gat), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT50), .B(new_n440_), .C1(new_n668_), .C2(new_n285_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(G1335gat));
  NAND4_X1  g491(.A1(new_n424_), .A2(new_n585_), .A3(new_n556_), .A4(new_n637_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT112), .Z(new_n694_));
  AOI21_X1  g493(.A(G85gat), .B1(new_n694_), .B2(new_n420_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n628_), .B1(new_n621_), .B2(KEYINPUT104), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n697_), .B(KEYINPUT43), .C1(new_n424_), .C2(new_n616_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n696_), .A2(new_n698_), .A3(new_n625_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(new_n671_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(new_n420_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n695_), .B1(new_n701_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g501(.A(G92gat), .B1(new_n694_), .B2(new_n362_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n422_), .A2(new_n345_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n700_), .B2(new_n704_), .ZN(G1337gat));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n381_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G99gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n694_), .A2(new_n381_), .A3(new_n480_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT114), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT51), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT114), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n707_), .A2(new_n714_), .A3(new_n708_), .A4(new_n709_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n711_), .A2(new_n713_), .A3(new_n715_), .ZN(G1338gat));
  NAND3_X1  g515(.A1(new_n694_), .A2(new_n475_), .A3(new_n285_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n699_), .A2(new_n285_), .A3(new_n671_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G106gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G106gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(G1339gat));
  INV_X1    g523(.A(KEYINPUT56), .ZN(new_n725_));
  INV_X1    g524(.A(new_n579_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n506_), .A2(new_n451_), .A3(new_n559_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n563_), .B1(new_n506_), .B2(new_n451_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n567_), .B1(new_n729_), .B2(new_n566_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n570_), .A2(KEYINPUT55), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n566_), .A2(new_n567_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT70), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n566_), .A2(KEYINPUT70), .A3(new_n567_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT55), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n729_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n730_), .B1(new_n731_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n726_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AOI211_X1 g540(.A(KEYINPUT117), .B(new_n730_), .C1(new_n731_), .C2(new_n738_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n725_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n729_), .A2(new_n566_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n572_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n570_), .A2(KEYINPUT55), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n737_), .B1(new_n736_), .B2(new_n729_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n745_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT117), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n739_), .A2(new_n740_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(KEYINPUT56), .A4(new_n726_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n743_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n581_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n554_), .A2(new_n555_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(KEYINPUT118), .A3(new_n755_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n580_), .A2(new_n581_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n541_), .A2(new_n543_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n536_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n545_), .A2(new_n538_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n762_), .B(new_n550_), .C1(new_n536_), .C2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n551_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n760_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT119), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n758_), .A2(new_n759_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n528_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT120), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n753_), .A2(new_n551_), .A3(new_n764_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n752_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT58), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n752_), .A2(KEYINPUT58), .A3(new_n773_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n616_), .A3(new_n777_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n769_), .A2(new_n770_), .B1(new_n771_), .B2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT58), .B1(new_n752_), .B2(new_n773_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n775_), .B(new_n772_), .C1(new_n743_), .C2(new_n751_), .ZN(new_n781_));
  NOR4_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n771_), .A4(new_n534_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n528_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT118), .B1(new_n752_), .B2(new_n755_), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n757_), .B(new_n754_), .C1(new_n743_), .C2(new_n751_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n786_), .B2(new_n767_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n782_), .B1(new_n787_), .B2(KEYINPUT57), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n472_), .B1(new_n779_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  INV_X1    g589(.A(new_n666_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n592_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n666_), .A2(KEYINPUT116), .A3(new_n584_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n534_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT121), .B1(new_n789_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n778_), .A2(new_n771_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n787_), .B2(KEYINPUT57), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n768_), .A2(KEYINPUT57), .A3(new_n528_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n776_), .A2(new_n616_), .A3(KEYINPUT120), .A4(new_n777_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n471_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804_));
  INV_X1    g603(.A(new_n796_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n285_), .A2(new_n401_), .A3(new_n362_), .A4(new_n380_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n797_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n557_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n800_), .A2(new_n778_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n787_), .A2(KEYINPUT57), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n471_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT122), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n814_), .B(new_n471_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n805_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n807_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n808_), .B2(new_n817_), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n809_), .B1(new_n821_), .B2(new_n557_), .ZN(G1340gat));
  OAI21_X1  g621(.A(G120gat), .B1(new_n819_), .B2(new_n586_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G120gat), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n797_), .A2(new_n806_), .A3(new_n807_), .A4(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G120gat), .B1(new_n592_), .B2(new_n824_), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n826_), .A2(KEYINPUT123), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT123), .B1(new_n826_), .B2(new_n827_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n823_), .A2(new_n830_), .ZN(G1341gat));
  AOI21_X1  g630(.A(G127gat), .B1(new_n808_), .B2(new_n472_), .ZN(new_n832_));
  INV_X1    g631(.A(G127gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n819_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n834_), .B2(new_n472_), .ZN(G1342gat));
  AOI21_X1  g634(.A(G134gat), .B1(new_n808_), .B2(new_n783_), .ZN(new_n836_));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n819_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n838_), .B2(new_n616_), .ZN(G1343gat));
  NAND4_X1  g638(.A1(new_n797_), .A2(new_n285_), .A3(new_n380_), .A4(new_n806_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n840_), .A2(new_n401_), .A3(new_n362_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n557_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G141gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n221_), .A3(new_n557_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n585_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT124), .B(G148gat), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n841_), .A2(new_n585_), .A3(new_n847_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1345gat));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n841_), .A2(new_n472_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n841_), .B2(new_n472_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1346gat));
  NAND2_X1  g654(.A1(new_n841_), .A2(new_n783_), .ZN(new_n856_));
  NOR4_X1   g655(.A1(new_n840_), .A2(new_n215_), .A3(new_n401_), .A4(new_n362_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n856_), .A2(new_n215_), .B1(new_n857_), .B2(new_n616_), .ZN(G1347gat));
  NOR2_X1   g657(.A1(new_n422_), .A2(new_n402_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n816_), .A2(new_n419_), .A3(new_n557_), .A4(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT62), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(G169gat), .A3(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n861_), .A2(KEYINPUT62), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n816_), .A2(new_n419_), .A3(new_n859_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n289_), .A3(new_n557_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n864_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n860_), .A2(G169gat), .A3(new_n869_), .A4(new_n862_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n865_), .A2(new_n868_), .A3(new_n870_), .ZN(G1348gat));
  AOI21_X1  g670(.A(G176gat), .B1(new_n867_), .B2(new_n592_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n797_), .A2(new_n806_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n873_), .A2(new_n290_), .A3(new_n285_), .A4(new_n586_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n859_), .B2(new_n874_), .ZN(G1349gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n285_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n422_), .A2(new_n402_), .A3(new_n471_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G183gat), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n866_), .A2(new_n471_), .A3(new_n307_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1350gat));
  OAI21_X1  g679(.A(G190gat), .B1(new_n866_), .B2(new_n534_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n783_), .A2(new_n308_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n866_), .B2(new_n882_), .ZN(G1351gat));
  AND2_X1   g682(.A1(new_n421_), .A2(new_n362_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n797_), .A2(new_n380_), .A3(new_n806_), .A4(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n556_), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n886_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n586_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g688(.A1(new_n885_), .A2(new_n471_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n890_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT63), .B(G211gat), .Z(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n890_), .B2(new_n892_), .ZN(G1354gat));
  AND3_X1   g692(.A1(new_n797_), .A2(new_n380_), .A3(new_n806_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n783_), .A4(new_n884_), .ZN(new_n896_));
  INV_X1    g695(.A(G218gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT126), .B1(new_n885_), .B2(new_n528_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n534_), .A2(new_n897_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT127), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n894_), .A2(new_n884_), .A3(new_n901_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n899_), .A2(new_n902_), .ZN(G1355gat));
endmodule


