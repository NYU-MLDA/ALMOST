//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  XOR2_X1   g000(.A(G127gat), .B(G155gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT16), .ZN(new_n203_));
  XOR2_X1   g002(.A(G183gat), .B(G211gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT17), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G57gat), .B(G64gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n209_));
  XOR2_X1   g008(.A(G71gat), .B(G78gat), .Z(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n210_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G231gat), .A2(G233gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n214_), .B(new_n215_), .Z(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT70), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218_));
  INV_X1    g017(.A(G1gat), .ZN(new_n219_));
  INV_X1    g018(.A(G8gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G1gat), .B(G8gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n217_), .B(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n225_), .A2(KEYINPUT17), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n207_), .B1(new_n226_), .B2(new_n205_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n225_), .A2(KEYINPUT71), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT12), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n214_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT7), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G106gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT6), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G99gat), .A2(G106gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT6), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n234_), .B(new_n238_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G85gat), .B(G92gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n246_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n238_), .A2(new_n234_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n241_), .B(KEYINPUT6), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n244_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n253_), .B(new_n254_), .C1(new_n258_), .C2(new_n250_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n245_), .A2(KEYINPUT9), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT10), .B(G99gat), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n237_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT64), .B(G92gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT9), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(G85gat), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n261_), .A2(new_n263_), .A3(new_n257_), .A4(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n233_), .B1(new_n260_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  AOI211_X1 g068(.A(KEYINPUT67), .B(new_n269_), .C1(new_n252_), .C2(new_n259_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n232_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n240_), .A2(new_n242_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n245_), .B1(new_n272_), .B2(new_n255_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n250_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n269_), .B1(new_n275_), .B2(new_n253_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n230_), .B1(new_n276_), .B2(new_n214_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n214_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(G230gat), .A2(G233gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n271_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n276_), .A2(new_n214_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n280_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT5), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G176gat), .B(G204gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n282_), .A2(new_n284_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n293_), .A2(KEYINPUT13), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(KEYINPUT13), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G190gat), .B(G218gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G134gat), .B(G162gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT36), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G232gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT34), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT35), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G29gat), .B(G36gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G43gat), .B(G50gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT15), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n259_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n254_), .B1(new_n275_), .B2(new_n253_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n267_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT67), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n260_), .A2(new_n233_), .A3(new_n267_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n312_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n276_), .A2(new_n310_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT68), .B1(new_n305_), .B2(new_n306_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n307_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n311_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n307_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n302_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n300_), .A2(KEYINPUT36), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n322_), .A2(new_n325_), .A3(KEYINPUT69), .A4(new_n327_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n326_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(KEYINPUT37), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT37), .ZN(new_n334_));
  AOI211_X1 g133(.A(new_n334_), .B(new_n326_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n229_), .A2(new_n297_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT72), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n311_), .A2(new_n224_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n310_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n224_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G229gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT73), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n224_), .B(new_n341_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(G229gat), .A3(G233gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G141gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G169gat), .B(G197gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  OR2_X1    g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n345_), .A2(new_n347_), .A3(new_n351_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G197gat), .A2(G204gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT21), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n361_));
  INV_X1    g160(.A(G211gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT81), .B1(new_n362_), .B2(G218gat), .ZN(new_n363_));
  INV_X1    g162(.A(G218gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(G211gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n359_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n358_), .B(KEYINPUT21), .C1(new_n365_), .C2(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT78), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G141gat), .A2(G148gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT2), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(G141gat), .A3(G148gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n381_), .A2(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n374_), .B1(new_n379_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n372_), .B1(KEYINPUT1), .B2(new_n370_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n370_), .A2(KEYINPUT1), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n380_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(new_n385_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n387_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n369_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n397_), .B(KEYINPUT80), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G78gat), .B(G106gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n369_), .B(new_n398_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT79), .B(KEYINPUT28), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n394_), .A2(new_n395_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G22gat), .B(G50gat), .Z(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n387_), .A2(new_n393_), .A3(KEYINPUT29), .ZN(new_n410_));
  INV_X1    g209(.A(new_n408_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n406_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n408_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n411_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n405_), .A3(new_n415_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(KEYINPUT83), .A2(new_n404_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n404_), .A2(KEYINPUT83), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n400_), .A2(new_n403_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n401_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT82), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n422_), .A3(new_n401_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n417_), .A2(new_n418_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n404_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G8gat), .B(G36gat), .Z(new_n428_));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT32), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G183gat), .A2(G190gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT23), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT23), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(G183gat), .A3(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G169gat), .A2(G176gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G176gat), .ZN(new_n445_));
  INV_X1    g244(.A(G169gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(KEYINPUT22), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT75), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n445_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT22), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G169gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(KEYINPUT22), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT75), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G183gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT25), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT25), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G183gat), .ZN(new_n458_));
  INV_X1    g257(.A(G190gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT26), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT26), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G190gat), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n456_), .A2(new_n458_), .A3(new_n460_), .A4(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(KEYINPUT24), .A3(new_n443_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT24), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n438_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT74), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n436_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n435_), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI22_X1  g273(.A1(new_n444_), .A2(new_n454_), .B1(new_n469_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT76), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n369_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT25), .B(G183gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT26), .B(G190gat), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n479_), .A2(new_n480_), .B1(new_n467_), .B2(new_n464_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n435_), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT74), .B1(new_n435_), .B2(KEYINPUT23), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n438_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n484_), .A3(new_n466_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n443_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n451_), .A2(KEYINPUT75), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT22), .B(G169gat), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n445_), .B(new_n488_), .C1(new_n489_), .C2(KEYINPUT75), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n485_), .A2(new_n491_), .A3(KEYINPUT76), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n477_), .A2(new_n478_), .A3(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G226gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n486_), .B1(new_n489_), .B2(new_n445_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(new_n474_), .B2(new_n440_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n481_), .A2(new_n466_), .A3(new_n439_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n498_), .B1(new_n502_), .B2(new_n369_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n493_), .A2(new_n497_), .A3(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n485_), .A2(KEYINPUT76), .A3(new_n491_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT76), .B1(new_n485_), .B2(new_n491_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n369_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n451_), .A2(new_n452_), .A3(new_n445_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n443_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n484_), .B2(new_n441_), .ZN(new_n511_));
  AND4_X1   g310(.A1(new_n466_), .A2(new_n463_), .A3(new_n468_), .A4(new_n439_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n508_), .B1(new_n513_), .B2(new_n478_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n497_), .B1(new_n507_), .B2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n434_), .B1(new_n504_), .B2(new_n515_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n505_), .A2(new_n506_), .A3(new_n369_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT20), .B1(new_n513_), .B2(new_n478_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n496_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(new_n478_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n496_), .A2(new_n498_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n507_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n522_), .A3(new_n433_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G127gat), .B(G134gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G113gat), .B(G120gat), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G113gat), .B(G120gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n387_), .B2(new_n393_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n381_), .A2(new_n383_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n385_), .A2(new_n384_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n376_), .A2(new_n378_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n373_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n528_), .A2(new_n530_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n390_), .A2(new_n392_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(KEYINPUT4), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G225gat), .A2(G233gat), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n538_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT4), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G1gat), .B(G29gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G85gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n532_), .A2(new_n542_), .A3(new_n540_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n547_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n547_), .B2(new_n554_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT90), .B1(new_n524_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n547_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n516_), .A4(new_n523_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n519_), .A2(new_n432_), .A3(new_n522_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n432_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n497_), .B1(new_n493_), .B2(new_n503_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n521_), .B1(new_n502_), .B2(new_n369_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n477_), .A2(new_n492_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(new_n369_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n568_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n547_), .A2(KEYINPUT33), .A3(new_n553_), .A4(new_n554_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n566_), .A2(new_n567_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT87), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n544_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n532_), .A2(KEYINPUT87), .A3(new_n540_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n543_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(KEYINPUT88), .A3(new_n552_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n552_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT88), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n541_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n575_), .B1(new_n581_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n427_), .B1(new_n564_), .B2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n561_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n568_), .B1(new_n504_), .B2(new_n515_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n590_), .A2(KEYINPUT27), .A3(new_n567_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT27), .B1(new_n567_), .B2(new_n573_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT30), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G71gat), .B(G99gat), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n597_), .A2(G43gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(G43gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n596_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n598_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n601_));
  OAI22_X1  g400(.A1(new_n505_), .A2(new_n506_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n600_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n477_), .A2(new_n603_), .A3(new_n492_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G227gat), .A2(G233gat), .ZN(new_n606_));
  INV_X1    g405(.A(G15gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT31), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n602_), .A2(new_n604_), .A3(new_n608_), .ZN(new_n612_));
  AND4_X1   g411(.A1(KEYINPUT77), .A2(new_n610_), .A3(new_n611_), .A4(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT77), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n611_), .B1(new_n615_), .B2(new_n612_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n538_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n610_), .A2(KEYINPUT77), .A3(new_n612_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT31), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n615_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n531_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n595_), .A2(new_n622_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n617_), .A2(new_n557_), .A3(new_n621_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT91), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n590_), .A2(KEYINPUT27), .A3(new_n567_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n567_), .A2(new_n573_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT91), .B(new_n627_), .C1(new_n628_), .C2(KEYINPUT27), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n624_), .A2(new_n630_), .A3(new_n427_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n354_), .B1(new_n623_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n338_), .A2(KEYINPUT72), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n339_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n219_), .A3(new_n561_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT38), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n296_), .A2(KEYINPUT92), .A3(new_n354_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT92), .B1(new_n296_), .B2(new_n354_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n229_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n330_), .A2(new_n331_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n326_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT93), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n584_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n628_), .A2(new_n644_), .A3(new_n574_), .A4(new_n566_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n646_), .A2(new_n427_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n622_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n631_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n643_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n639_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n219_), .B1(new_n651_), .B2(new_n561_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT94), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n636_), .A2(new_n653_), .ZN(G1324gat));
  INV_X1    g453(.A(new_n630_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G8gat), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n657_), .A2(new_n658_), .A3(KEYINPUT39), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT95), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(new_n662_), .A3(KEYINPUT39), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n657_), .B2(KEYINPUT39), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n659_), .A2(new_n661_), .A3(new_n663_), .A4(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n634_), .A2(new_n220_), .A3(new_n655_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n667_), .B(new_n669_), .ZN(G1325gat));
  AOI21_X1  g469(.A(new_n607_), .B1(new_n651_), .B2(new_n648_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT41), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n634_), .A2(new_n607_), .A3(new_n648_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(G22gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n427_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n651_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT99), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT98), .B(KEYINPUT42), .Z(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n634_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1327gat));
  XOR2_X1   g481(.A(new_n227_), .B(new_n228_), .Z(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n332_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(new_n296_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n632_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(G29gat), .A3(new_n557_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n648_), .B1(new_n588_), .B2(new_n594_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n624_), .A2(new_n630_), .A3(new_n427_), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n689_), .A2(new_n690_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT100), .B(KEYINPUT43), .Z(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT101), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n691_), .A2(new_n696_), .A3(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n642_), .A2(new_n334_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n332_), .A2(KEYINPUT37), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n649_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n700_), .A2(new_n649_), .A3(KEYINPUT102), .A4(new_n701_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n695_), .A2(new_n697_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n637_), .A2(new_n683_), .A3(new_n638_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n688_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n623_), .A2(new_n631_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT102), .B1(new_n710_), .B2(new_n701_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n705_), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT101), .B(new_n692_), .C1(new_n700_), .C2(new_n649_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n696_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n714_));
  OAI22_X1  g513(.A1(new_n711_), .A2(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n707_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(KEYINPUT103), .A3(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n708_), .A2(new_n709_), .A3(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(KEYINPUT44), .A3(new_n716_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n561_), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n687_), .B1(new_n720_), .B2(G29gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT104), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n718_), .A2(new_n655_), .A3(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n686_), .A2(G36gat), .A3(new_n630_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT46), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT105), .B(new_n731_), .C1(new_n724_), .C2(new_n727_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1329gat));
  XNOR2_X1  g532(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G43gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n622_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n718_), .A2(new_n719_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n736_), .B1(new_n686_), .B2(new_n622_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n735_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n738_), .A2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT107), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n734_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n743_), .A2(new_n747_), .ZN(G1330gat));
  OR3_X1    g547(.A1(new_n686_), .A2(G50gat), .A3(new_n427_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n718_), .A2(new_n676_), .A3(new_n719_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n750_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT108), .B1(new_n750_), .B2(G50gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n751_), .B2(new_n752_), .ZN(G1331gat));
  INV_X1    g552(.A(new_n354_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n297_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n649_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n756_), .A2(new_n683_), .A3(new_n700_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT109), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT109), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n561_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(G57gat), .ZN(new_n761_));
  NOR4_X1   g560(.A1(new_n650_), .A2(new_n683_), .A3(new_n754_), .A4(new_n297_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n557_), .A2(new_n761_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n760_), .A2(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(G1332gat));
  INV_X1    g563(.A(G64gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n762_), .B2(new_n655_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT48), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n757_), .A2(new_n765_), .A3(new_n655_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1333gat));
  INV_X1    g568(.A(G71gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n762_), .B2(new_n648_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT49), .Z(new_n772_));
  NAND3_X1  g571(.A1(new_n757_), .A2(new_n770_), .A3(new_n648_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1334gat));
  INV_X1    g573(.A(G78gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n762_), .B2(new_n676_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT50), .Z(new_n777_));
  NAND3_X1  g576(.A1(new_n757_), .A2(new_n775_), .A3(new_n676_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1335gat));
  OR2_X1    g578(.A1(new_n684_), .A2(new_n756_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT110), .ZN(new_n781_));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n561_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n683_), .A2(new_n755_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n695_), .A2(new_n697_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n704_), .A2(new_n705_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n561_), .A2(G85gat), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT111), .Z(new_n788_));
  AOI21_X1  g587(.A(new_n782_), .B1(new_n786_), .B2(new_n788_), .ZN(G1336gat));
  AOI21_X1  g588(.A(G92gat), .B1(new_n781_), .B2(new_n655_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n655_), .A2(new_n264_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n786_), .B2(new_n791_), .ZN(G1337gat));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n648_), .A3(new_n262_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n706_), .A2(new_n622_), .A3(new_n783_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n236_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT51), .ZN(G1338gat));
  AND3_X1   g595(.A1(new_n781_), .A2(new_n237_), .A3(new_n676_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n237_), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n786_), .B2(new_n676_), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n706_), .A2(KEYINPUT112), .A3(new_n427_), .A4(new_n783_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n798_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n803_), .B(new_n798_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n797_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n808_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n810_), .B(new_n797_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n338_), .A2(new_n813_), .A3(new_n354_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT54), .B1(new_n337_), .B2(new_n754_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n351_), .B1(new_n346_), .B2(new_n344_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n344_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n340_), .A2(new_n342_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n353_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n353_), .A2(new_n822_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT116), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n293_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n282_), .A2(KEYINPUT55), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n271_), .A2(new_n281_), .A3(new_n829_), .A4(new_n277_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n271_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n280_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n289_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(KEYINPUT115), .A3(new_n836_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n828_), .A2(new_n830_), .B1(new_n280_), .B2(new_n832_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n835_), .B1(new_n838_), .B2(new_n289_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  INV_X1    g639(.A(new_n836_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n838_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n837_), .A2(new_n839_), .A3(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n354_), .A2(new_n291_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n827_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n818_), .B1(new_n845_), .B2(new_n332_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT117), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n848_), .B(new_n818_), .C1(new_n845_), .C2(new_n332_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n843_), .A2(new_n844_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT57), .B(new_n642_), .C1(new_n851_), .C2(new_n827_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n826_), .A2(new_n824_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n290_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n853_), .B2(new_n290_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n839_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n838_), .A2(new_n841_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT58), .B(new_n857_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n700_), .A3(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n852_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n850_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n229_), .B1(new_n866_), .B2(KEYINPUT119), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n852_), .A2(new_n864_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n817_), .B1(new_n867_), .B2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n655_), .A2(new_n676_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n622_), .A2(new_n557_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G113gat), .B1(new_n876_), .B2(new_n754_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n852_), .A2(new_n864_), .A3(new_n846_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n879_), .A2(KEYINPUT120), .A3(new_n683_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT120), .B1(new_n879_), .B2(new_n683_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n817_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n875_), .A2(KEYINPUT59), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n878_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n879_), .A2(new_n683_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n816_), .B1(new_n886_), .B2(KEYINPUT120), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT121), .B(new_n883_), .C1(new_n887_), .C2(new_n880_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT59), .B1(new_n872_), .B2(new_n875_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(G113gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n754_), .B2(KEYINPUT122), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(KEYINPUT122), .B2(new_n892_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n877_), .B1(new_n891_), .B2(new_n894_), .ZN(G1340gat));
  NAND3_X1  g694(.A1(new_n889_), .A2(new_n296_), .A3(new_n890_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G120gat), .ZN(new_n897_));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n297_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n876_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n897_), .A2(new_n900_), .ZN(G1341gat));
  NAND3_X1  g700(.A1(new_n889_), .A2(new_n229_), .A3(new_n890_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G127gat), .ZN(new_n903_));
  INV_X1    g702(.A(new_n876_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n904_), .A2(G127gat), .A3(new_n683_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1342gat));
  NAND3_X1  g705(.A1(new_n889_), .A2(new_n700_), .A3(new_n890_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G134gat), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n904_), .A2(G134gat), .A3(new_n643_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1343gat));
  NOR4_X1   g709(.A1(new_n655_), .A2(new_n648_), .A3(new_n557_), .A4(new_n427_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n872_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n754_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n296_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT123), .B(G148gat), .Z(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1345gat));
  NAND2_X1  g717(.A1(new_n913_), .A2(new_n229_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT61), .B(G155gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1346gat));
  INV_X1    g720(.A(G162gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n913_), .B2(new_n700_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n683_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n866_), .A2(KEYINPUT119), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n816_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n643_), .A2(G162gat), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n926_), .A2(new_n911_), .A3(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT124), .B1(new_n923_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n928_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n926_), .A2(new_n911_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G162gat), .B1(new_n931_), .B2(new_n336_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n930_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n929_), .A2(new_n934_), .ZN(G1347gat));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n655_), .A2(new_n427_), .A3(new_n624_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n882_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n754_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n936_), .B1(new_n939_), .B2(G169gat), .ZN(new_n940_));
  AOI211_X1 g739(.A(KEYINPUT62), .B(new_n446_), .C1(new_n938_), .C2(new_n754_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n938_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n754_), .A2(new_n489_), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n943_), .B(KEYINPUT125), .Z(new_n944_));
  OAI22_X1  g743(.A1(new_n940_), .A2(new_n941_), .B1(new_n942_), .B2(new_n944_), .ZN(G1348gat));
  AOI21_X1  g744(.A(G176gat), .B1(new_n938_), .B2(new_n296_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n872_), .A2(new_n937_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n297_), .A2(new_n445_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n946_), .B1(new_n947_), .B2(new_n948_), .ZN(G1349gat));
  AOI21_X1  g748(.A(G183gat), .B1(new_n947_), .B2(new_n229_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n683_), .A2(new_n479_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n938_), .B2(new_n951_), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n942_), .B2(new_n336_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n480_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n643_), .A2(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n953_), .B1(new_n942_), .B2(new_n955_), .ZN(G1351gat));
  NAND3_X1  g755(.A1(new_n655_), .A2(new_n589_), .A3(new_n622_), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT126), .B1(new_n872_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959_));
  INV_X1    g758(.A(new_n957_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n926_), .A2(new_n959_), .A3(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n958_), .A2(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(G197gat), .B1(new_n962_), .B2(new_n754_), .ZN(new_n963_));
  INV_X1    g762(.A(G197gat), .ZN(new_n964_));
  AOI211_X1 g763(.A(new_n964_), .B(new_n354_), .C1(new_n958_), .C2(new_n961_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n963_), .A2(new_n965_), .ZN(G1352gat));
  NOR3_X1   g765(.A1(new_n872_), .A2(KEYINPUT126), .A3(new_n957_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n959_), .B1(new_n926_), .B2(new_n960_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n296_), .B1(new_n967_), .B2(new_n968_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(KEYINPUT127), .B(G204gat), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n969_), .A2(new_n971_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n962_), .A2(new_n296_), .A3(new_n970_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(G1353gat));
  OR2_X1    g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n975_), .B1(new_n962_), .B2(new_n229_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(KEYINPUT63), .B(G211gat), .ZN(new_n977_));
  AOI211_X1 g776(.A(new_n683_), .B(new_n977_), .C1(new_n958_), .C2(new_n961_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n976_), .A2(new_n978_), .ZN(G1354gat));
  NOR2_X1   g778(.A1(new_n643_), .A2(G218gat), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n962_), .A2(new_n980_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n336_), .B1(new_n958_), .B2(new_n961_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n364_), .B2(new_n982_), .ZN(G1355gat));
endmodule


