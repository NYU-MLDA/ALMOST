//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT104), .ZN(new_n203_));
  OR2_X1    g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G218gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G211gat), .ZN(new_n210_));
  INV_X1    g009(.A(G211gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G218gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT90), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(new_n212_), .A3(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n208_), .A2(new_n214_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n217_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n216_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n215_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT92), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT92), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n218_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(G176gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT24), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT95), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  INV_X1    g037(.A(G183gat), .ZN(new_n239_));
  INV_X1    g038(.A(G190gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n229_), .A2(KEYINPUT95), .A3(new_n234_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n237_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n239_), .A2(new_n240_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n241_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G169gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n233_), .C1(new_n252_), .C2(G176gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n224_), .A2(new_n226_), .A3(new_n248_), .A4(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n223_), .A2(KEYINPUT91), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT79), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G183gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n257_), .A2(KEYINPUT25), .B1(new_n258_), .B2(G190gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT80), .B1(new_n258_), .B2(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n240_), .A3(KEYINPUT26), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n259_), .B(new_n263_), .C1(KEYINPUT25), .C2(new_n257_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT81), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n245_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n241_), .A2(new_n244_), .A3(KEYINPUT81), .A4(new_n242_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n264_), .A2(new_n234_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n250_), .A2(KEYINPUT83), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT82), .B(G169gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT22), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n231_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n241_), .A2(new_n274_), .A3(new_n242_), .A4(new_n249_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n270_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n269_), .A2(new_n273_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n268_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT91), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n218_), .A2(new_n222_), .A3(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n255_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n254_), .A2(new_n281_), .A3(KEYINPUT20), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT102), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT19), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT20), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n248_), .A2(new_n253_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n223_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n280_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n279_), .B1(new_n218_), .B2(new_n222_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n268_), .B(new_n277_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n285_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n289_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n283_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n286_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT18), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n203_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n282_), .A2(new_n285_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(new_n294_), .A3(KEYINPUT102), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n304_), .A2(new_n203_), .A3(new_n301_), .A4(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT27), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n248_), .A2(new_n218_), .A3(new_n222_), .A4(new_n253_), .ZN(new_n308_));
  AND4_X1   g107(.A1(KEYINPUT20), .A2(new_n281_), .A3(new_n293_), .A4(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n293_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n307_), .B1(new_n311_), .B2(new_n300_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n202_), .B1(new_n302_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n304_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT104), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n316_), .A2(KEYINPUT105), .A3(new_n306_), .A4(new_n312_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n311_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n301_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n311_), .A2(new_n300_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n314_), .A2(new_n317_), .B1(new_n307_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT97), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OR3_X1    g126(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT88), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n331_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n327_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OR3_X1    g135(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n337_), .A2(new_n338_), .B1(G141gat), .B2(G148gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n324_), .B1(new_n326_), .B2(KEYINPUT1), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(KEYINPUT1), .B2(new_n324_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT87), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT87), .B1(new_n339_), .B2(new_n341_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n336_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT89), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT89), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n346_), .B(new_n336_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G127gat), .B(G134gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n347_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n339_), .A2(new_n341_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT87), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT87), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n334_), .A2(new_n335_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n355_), .A2(new_n356_), .B1(new_n357_), .B2(new_n327_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n350_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n345_), .A2(new_n347_), .A3(new_n351_), .A4(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n323_), .B1(new_n361_), .B2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n360_), .A2(KEYINPUT97), .A3(new_n365_), .A4(new_n363_), .ZN(new_n368_));
  XOR2_X1   g167(.A(KEYINPUT98), .B(KEYINPUT0), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT99), .ZN(new_n370_));
  XOR2_X1   g169(.A(G1gat), .B(G29gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G57gat), .B(G85gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  NAND3_X1  g173(.A1(new_n352_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n367_), .A2(new_n368_), .A3(new_n374_), .A4(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT103), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n368_), .A2(new_n375_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT103), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n374_), .A4(new_n367_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n374_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n367_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(new_n378_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n377_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n345_), .A2(new_n347_), .A3(KEYINPUT29), .ZN(new_n387_));
  AND2_X1   g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n290_), .A2(new_n388_), .A3(new_n291_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n344_), .A2(KEYINPUT29), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n224_), .A2(new_n226_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n387_), .A2(new_n389_), .B1(new_n392_), .B2(new_n388_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n386_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n345_), .B2(new_n347_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G22gat), .B(G50gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT28), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n397_), .B(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT94), .B1(new_n396_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n387_), .A2(new_n389_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n392_), .A2(new_n388_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n395_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT93), .ZN(new_n405_));
  INV_X1    g204(.A(new_n399_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n397_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT94), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n393_), .B(new_n394_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n401_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n401_), .B2(new_n409_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n322_), .A2(new_n385_), .A3(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n352_), .A2(KEYINPUT101), .A3(new_n359_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT101), .B1(new_n352_), .B2(new_n359_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n364_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n360_), .A2(new_n364_), .A3(new_n363_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n382_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n319_), .B(new_n320_), .C1(new_n417_), .C2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT100), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n376_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n422_), .B2(KEYINPUT33), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n376_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n377_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n300_), .A2(KEYINPUT32), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n318_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n427_), .B2(new_n296_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n423_), .A2(new_n425_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n414_), .B1(new_n430_), .B2(new_n413_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n278_), .B(KEYINPUT85), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT31), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT84), .B1(new_n350_), .B2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n433_), .B2(new_n350_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G71gat), .B(G99gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G43gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n435_), .B(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G227gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(G15gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT30), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n438_), .A2(new_n442_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n432_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n438_), .A2(new_n442_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n432_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n438_), .A2(new_n442_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n411_), .A2(new_n412_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n314_), .A2(new_n317_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n321_), .A2(new_n307_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n385_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT106), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT106), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n322_), .A2(new_n456_), .A3(new_n451_), .A4(new_n385_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n431_), .A2(new_n450_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G1gat), .A2(G8gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT14), .ZN(new_n461_));
  INV_X1    g260(.A(G22gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n440_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G15gat), .A2(G22gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G1gat), .ZN(new_n466_));
  INV_X1    g265(.A(G8gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT76), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n460_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n468_), .B2(new_n460_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n461_), .B(new_n465_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n472_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n465_), .A2(new_n461_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n459_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G29gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n481_), .A2(KEYINPUT15), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT15), .B1(new_n481_), .B2(new_n482_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n473_), .A2(new_n476_), .A3(new_n459_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n478_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n481_), .A2(new_n482_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n486_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(new_n477_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT78), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT78), .ZN(new_n495_));
  INV_X1    g294(.A(new_n488_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n478_), .A2(new_n496_), .A3(new_n486_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n492_), .B1(new_n490_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n493_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n493_), .B(new_n504_), .C1(new_n495_), .C2(new_n498_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G230gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT64), .ZN(new_n510_));
  INV_X1    g309(.A(G99gat), .ZN(new_n511_));
  INV_X1    g310(.A(G106gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT7), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(KEYINPUT64), .A2(G99gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n512_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n514_), .A2(new_n519_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G85gat), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT65), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(KEYINPUT66), .B2(KEYINPUT8), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n530_), .B2(KEYINPUT8), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n523_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n512_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n526_), .A2(KEYINPUT9), .A3(new_n527_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n527_), .A2(KEYINPUT9), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n519_), .A2(new_n536_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n539_));
  NOR4_X1   g338(.A1(KEYINPUT64), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n521_), .B1(new_n520_), .B2(new_n512_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n528_), .B1(new_n542_), .B2(new_n519_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n531_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n533_), .B(new_n539_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT67), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n544_), .B1(new_n523_), .B2(new_n529_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n533_), .A4(new_n539_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G71gat), .B(G78gat), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT11), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(KEYINPUT11), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n551_), .A2(KEYINPUT11), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n553_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n546_), .A2(new_n550_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n509_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(KEYINPUT12), .B(new_n553_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n545_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT68), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT68), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n545_), .A2(new_n572_), .A3(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n574_), .B(new_n559_), .C1(KEYINPUT12), .C2(new_n561_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n562_), .B(new_n567_), .C1(new_n575_), .C2(new_n509_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT69), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n546_), .A2(new_n550_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n558_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT12), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n582_), .A2(new_n508_), .A3(new_n559_), .A4(new_n574_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n583_), .A2(KEYINPUT69), .A3(new_n562_), .A4(new_n567_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n562_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n566_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n585_), .A2(KEYINPUT13), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT13), .B1(new_n585_), .B2(new_n587_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n458_), .A2(new_n507_), .A3(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G190gat), .B(G218gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT73), .ZN(new_n594_));
  XOR2_X1   g393(.A(G134gat), .B(G162gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT36), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n546_), .A2(new_n488_), .A3(new_n550_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT72), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n485_), .A2(new_n545_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT72), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n546_), .A2(new_n601_), .A3(new_n550_), .A4(new_n488_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT34), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT35), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n599_), .A2(new_n600_), .A3(new_n602_), .A4(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n599_), .A2(KEYINPUT71), .A3(new_n602_), .A4(new_n605_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(KEYINPUT35), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT70), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n606_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n597_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n599_), .A2(new_n602_), .A3(new_n605_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n615_), .B(new_n600_), .C1(KEYINPUT71), .C2(new_n609_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n596_), .A4(new_n611_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n614_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n614_), .B2(new_n618_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n478_), .A2(new_n486_), .ZN(new_n623_));
  AND2_X1   g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n558_), .B(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(new_n630_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT17), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n623_), .A2(new_n625_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n626_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n634_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n626_), .B2(new_n635_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n622_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n592_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n466_), .A3(new_n426_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n614_), .A2(new_n618_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n642_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n592_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n385_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n645_), .A2(new_n646_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n647_), .A2(new_n652_), .A3(new_n653_), .ZN(G1324gat));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n467_), .B1(new_n655_), .B2(KEYINPUT39), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n656_), .B1(new_n651_), .B2(new_n322_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(KEYINPUT107), .A3(new_n658_), .ZN(new_n659_));
  OAI221_X1 g458(.A(new_n656_), .B1(new_n655_), .B2(KEYINPUT39), .C1(new_n651_), .C2(new_n322_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n322_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n644_), .A2(new_n467_), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(G1325gat));
  INV_X1    g464(.A(new_n450_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n644_), .A2(new_n440_), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n592_), .A2(new_n666_), .A3(new_n650_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT41), .B1(new_n668_), .B2(G15gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT108), .ZN(G1326gat));
  NAND3_X1  g471(.A1(new_n644_), .A2(new_n462_), .A3(new_n413_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n592_), .A2(new_n413_), .A3(new_n650_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(G22gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1327gat));
  NOR2_X1   g477(.A1(new_n648_), .A2(new_n641_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n592_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n426_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n621_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n614_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n458_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n455_), .A2(new_n457_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n426_), .A2(new_n429_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n422_), .A2(KEYINPUT33), .ZN(new_n689_));
  INV_X1    g488(.A(new_n420_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n425_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n413_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n666_), .B1(new_n694_), .B2(new_n414_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n686_), .B(new_n622_), .C1(new_n687_), .C2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n685_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n591_), .A2(new_n507_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n642_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n702_), .B(new_n699_), .C1(new_n685_), .C2(new_n696_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n426_), .A2(G29gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n681_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n704_), .B2(new_n661_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n592_), .A2(new_n708_), .A3(new_n661_), .A4(new_n679_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n712_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n701_), .A2(new_n703_), .A3(new_n322_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n714_), .B(KEYINPUT46), .C1(new_n708_), .C2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(G1329gat));
  NAND2_X1  g516(.A1(new_n666_), .A2(G43gat), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n701_), .A2(new_n703_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(G43gat), .B1(new_n680_), .B2(new_n666_), .ZN(new_n720_));
  OR3_X1    g519(.A1(new_n719_), .A2(KEYINPUT47), .A3(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT47), .B1(new_n719_), .B2(new_n720_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n680_), .B2(new_n413_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n413_), .A2(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n704_), .B2(new_n725_), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n591_), .A2(new_n507_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n458_), .A2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n650_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(G57gat), .A3(new_n426_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT110), .Z(new_n731_));
  AND2_X1   g530(.A1(new_n728_), .A2(new_n643_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n426_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1332gat));
  NOR2_X1   g533(.A1(new_n322_), .A2(G64gat), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT111), .Z(new_n736_));
  NAND2_X1  g535(.A1(new_n732_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n728_), .A2(new_n661_), .A3(new_n650_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G64gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT112), .Z(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n732_), .A2(new_n744_), .A3(new_n666_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n729_), .A2(new_n666_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G71gat), .ZN(new_n747_));
  XOR2_X1   g546(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(new_n748_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n745_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n732_), .A2(new_n752_), .A3(new_n413_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n729_), .A2(new_n413_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G78gat), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n755_), .A2(new_n756_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n728_), .A2(new_n760_), .A3(new_n679_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n728_), .B2(new_n679_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n524_), .A3(new_n426_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n591_), .A2(new_n507_), .A3(new_n642_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n685_), .B2(new_n696_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(new_n426_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n524_), .B2(new_n768_), .ZN(G1336gat));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n525_), .A3(new_n661_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n767_), .A2(new_n661_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n525_), .B2(new_n771_), .ZN(G1337gat));
  AND2_X1   g571(.A1(new_n534_), .A2(new_n535_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n764_), .A2(new_n773_), .A3(new_n666_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n767_), .A2(new_n666_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n511_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT51), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n764_), .A2(new_n773_), .A3(new_n666_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n778_), .B(new_n779_), .C1(new_n511_), .C2(new_n775_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1338gat));
  OAI211_X1 g580(.A(new_n512_), .B(new_n413_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  OAI21_X1  g582(.A(G106gat), .B1(new_n783_), .B2(KEYINPUT116), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n767_), .B2(new_n413_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(KEYINPUT116), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n786_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT53), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n785_), .A2(new_n786_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n788_), .A4(new_n782_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1339gat));
  NAND2_X1  g593(.A1(new_n585_), .A2(new_n506_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n573_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n572_), .B1(new_n545_), .B2(new_n569_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n559_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n798_), .A2(new_n581_), .A3(new_n509_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n509_), .B1(new_n798_), .B2(new_n581_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(KEYINPUT55), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n575_), .A2(new_n802_), .A3(new_n509_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n566_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n800_), .A2(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n583_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n799_), .A2(KEYINPUT55), .A3(new_n800_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n795_), .B1(new_n806_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n490_), .A2(new_n497_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n502_), .B1(new_n813_), .B2(new_n492_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT118), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n487_), .A2(new_n490_), .A3(G229gat), .A4(G233gat), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n814_), .A2(KEYINPUT118), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n503_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n648_), .B1(new_n812_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(new_n578_), .B2(new_n584_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n566_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n805_), .B(new_n567_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT58), .B(new_n824_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n622_), .A3(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT57), .B(new_n648_), .C1(new_n812_), .C2(new_n820_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n823_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n642_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n589_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n503_), .A2(new_n641_), .A3(new_n505_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT117), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n503_), .A2(new_n641_), .A3(new_n838_), .A4(new_n505_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n585_), .A2(KEYINPUT13), .A3(new_n587_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n835_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n843_), .A2(new_n622_), .A3(KEYINPUT54), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n588_), .A2(new_n589_), .A3(new_n840_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n684_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n385_), .B1(new_n834_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n322_), .A2(new_n451_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(KEYINPUT59), .A3(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n507_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n507_), .A2(G113gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n853_), .B2(new_n860_), .ZN(G1340gat));
  INV_X1    g660(.A(new_n853_), .ZN(new_n862_));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n590_), .B2(KEYINPUT60), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n862_), .B(new_n864_), .C1(KEYINPUT60), .C2(new_n863_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n590_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT119), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n865_), .B(new_n869_), .C1(new_n866_), .C2(new_n863_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1341gat));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n853_), .B2(new_n642_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(KEYINPUT120), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n873_), .A2(KEYINPUT120), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n642_), .A2(new_n872_), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n874_), .B(new_n875_), .C1(new_n857_), .C2(new_n876_), .ZN(G1342gat));
  OAI21_X1  g676(.A(G134gat), .B1(new_n858_), .B2(new_n684_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n648_), .A2(G134gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n853_), .B2(new_n879_), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n661_), .A2(new_n693_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n450_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n881_), .B1(new_n850_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n848_), .B1(new_n833_), .B2(new_n642_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n886_), .A2(KEYINPUT121), .A3(new_n385_), .A4(new_n883_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n506_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g688(.A(new_n591_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g690(.A(new_n641_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT122), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n894_), .B(new_n641_), .C1(new_n885_), .C2(new_n887_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n893_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1346gat));
  NOR2_X1   g698(.A1(new_n885_), .A2(new_n887_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G162gat), .B1(new_n900_), .B2(new_n684_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n648_), .A2(G162gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n900_), .B2(new_n902_), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n834_), .A2(new_n849_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n322_), .A2(new_n426_), .A3(new_n450_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n905_), .A2(KEYINPUT123), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(KEYINPUT123), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n413_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n909_), .A2(new_n507_), .A3(new_n252_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n909_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n230_), .B1(new_n911_), .B2(new_n506_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n912_), .B2(KEYINPUT62), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(KEYINPUT62), .B2(new_n912_), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n909_), .A2(new_n590_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n231_), .A2(KEYINPUT124), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n231_), .A2(KEYINPUT124), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n915_), .B2(new_n917_), .ZN(G1349gat));
  NOR2_X1   g718(.A1(new_n909_), .A2(new_n642_), .ZN(new_n920_));
  MUX2_X1   g719(.A(G183gat), .B(new_n227_), .S(new_n920_), .Z(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n909_), .B2(new_n684_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n649_), .A2(new_n228_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT125), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n909_), .B2(new_n924_), .ZN(G1351gat));
  NAND3_X1  g724(.A1(new_n413_), .A2(new_n385_), .A3(new_n450_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n886_), .A2(new_n322_), .A3(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n506_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n591_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g730(.A(new_n642_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n932_), .B(KEYINPUT126), .Z(new_n933_));
  NAND2_X1  g732(.A1(new_n927_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n934_), .B(new_n935_), .Z(G1354gat));
  NAND3_X1  g735(.A1(new_n927_), .A2(new_n209_), .A3(new_n649_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n927_), .A2(new_n622_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n209_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


