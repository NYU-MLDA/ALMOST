//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  NOR3_X1   g000(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT25), .B(G183gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G190gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT24), .A4(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n205_), .A2(new_n207_), .A3(new_n212_), .A4(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(new_n217_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT81), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n228_), .A2(new_n209_), .A3(G183gat), .A4(G190gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n224_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n219_), .A2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT82), .B(G15gat), .Z(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G127gat), .B(G134gat), .Z(new_n237_));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  XNOR2_X1  g038(.A(new_n236_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G71gat), .B(G99gat), .ZN(new_n241_));
  INV_X1    g040(.A(G43gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT30), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT31), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n240_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G8gat), .B(G36gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G64gat), .B(G92gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n254_), .A2(KEYINPUT32), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT19), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n225_), .A2(KEYINPUT25), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(G183gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n226_), .A2(KEYINPUT26), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT26), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(G190gat), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .A4(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n216_), .B(new_n213_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT91), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n224_), .A2(new_n229_), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n216_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT91), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n265_), .A2(new_n268_), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n212_), .A2(new_n207_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n227_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n223_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT21), .ZN(new_n281_));
  AND2_X1   g080(.A1(G197gat), .A2(G204gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G197gat), .A2(G204gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G197gat), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G197gat), .A2(G204gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT21), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n284_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G218gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G211gat), .ZN(new_n293_));
  INV_X1    g092(.A(G211gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G218gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(KEYINPUT21), .A3(new_n287_), .A4(new_n288_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n280_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT20), .ZN(new_n300_));
  INV_X1    g099(.A(new_n202_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n218_), .A2(new_n265_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n277_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n302_), .A2(new_n303_), .B1(new_n223_), .B2(new_n230_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n291_), .A2(new_n297_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n258_), .B1(new_n299_), .B2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n300_), .B1(new_n232_), .B2(new_n298_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n276_), .A2(new_n305_), .A3(new_n279_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n258_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n255_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n299_), .A2(new_n258_), .A3(new_n306_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n308_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n298_), .B1(new_n280_), .B2(KEYINPUT95), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n276_), .A2(new_n315_), .A3(new_n279_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n312_), .B1(new_n317_), .B2(new_n258_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n311_), .B1(new_n318_), .B2(new_n255_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G85gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT0), .B(G57gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G155gat), .B(G162gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(KEYINPUT1), .ZN(new_n326_));
  OR2_X1    g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT85), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n328_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT84), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n325_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n332_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n325_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n337_), .A2(new_n338_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n335_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n340_), .B(KEYINPUT84), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n346_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(KEYINPUT86), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n239_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n331_), .B1(new_n350_), .B2(KEYINPUT86), .ZN(new_n353_));
  INV_X1    g152(.A(new_n239_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n343_), .A2(new_n344_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n356_), .A3(KEYINPUT4), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n353_), .A2(new_n355_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n239_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n324_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n368_), .A2(new_n323_), .A3(new_n365_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n319_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n323_), .B(new_n371_), .C1(new_n368_), .C2(new_n365_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n253_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n305_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n305_), .A2(new_n219_), .A3(new_n231_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT20), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n257_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n308_), .A2(new_n309_), .A3(new_n258_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n254_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n352_), .A2(new_n356_), .A3(new_n363_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT94), .B1(new_n382_), .B2(new_n324_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT94), .A3(new_n324_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n384_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n372_), .B(new_n381_), .C1(new_n383_), .C2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n367_), .A2(new_n371_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n370_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n350_), .A2(KEYINPUT86), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(new_n355_), .A3(new_n391_), .A4(new_n332_), .ZN(new_n392_));
  XOR2_X1   g191(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G22gat), .B(G50gat), .Z(new_n395_));
  INV_X1    g194(.A(new_n393_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n353_), .A2(new_n391_), .A3(new_n355_), .A4(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n394_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n389_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n397_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n395_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n394_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT89), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n358_), .A2(KEYINPUT29), .ZN(new_n406_));
  OAI211_X1 g205(.A(G228gat), .B(G233gat), .C1(new_n305_), .C2(KEYINPUT88), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n298_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n391_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(new_n305_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n400_), .B(new_n405_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT89), .B1(new_n403_), .B2(new_n404_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n416_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n414_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n388_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT96), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n364_), .A2(new_n324_), .A3(new_n366_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n323_), .B1(new_n368_), .B2(new_n365_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(KEYINPUT96), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n417_), .A2(new_n420_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n379_), .A2(KEYINPUT27), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n318_), .B2(new_n253_), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n377_), .A2(new_n254_), .A3(new_n378_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n254_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT98), .B(new_n433_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n431_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n428_), .A2(new_n429_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n248_), .B1(new_n422_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n246_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT99), .B(new_n431_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT99), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n438_), .A2(new_n439_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n318_), .A2(new_n253_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n430_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n421_), .B(new_n443_), .C1(new_n444_), .C2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT100), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT98), .B1(new_n380_), .B2(new_n433_), .ZN(new_n454_));
  AOI211_X1 g253(.A(new_n437_), .B(new_n432_), .C1(new_n373_), .C2(new_n379_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n449_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT99), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n440_), .A2(new_n445_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n459_), .A2(KEYINPUT100), .A3(new_n421_), .A4(new_n443_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n442_), .B1(new_n453_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G29gat), .B(G36gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G43gat), .B(G50gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT15), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467_));
  INV_X1    g266(.A(G1gat), .ZN(new_n468_));
  INV_X1    g267(.A(G8gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G8gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n466_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n465_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G229gat), .A2(G233gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n473_), .B(new_n465_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n477_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT78), .ZN(new_n484_));
  XOR2_X1   g283(.A(G169gat), .B(G197gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n487_), .A2(KEYINPUT77), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n482_), .B(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n461_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G230gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT64), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT7), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT6), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G85gat), .B(G92gat), .Z(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT8), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(KEYINPUT65), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n493_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n504_), .A3(new_n496_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n498_), .A2(KEYINPUT8), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n499_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT10), .B(G99gat), .Z(new_n508_));
  INV_X1    g307(.A(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n498_), .A2(KEYINPUT9), .ZN(new_n511_));
  INV_X1    g310(.A(G85gat), .ZN(new_n512_));
  INV_X1    g311(.A(G92gat), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT9), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .A4(new_n496_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G57gat), .B(G64gat), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(KEYINPUT11), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(KEYINPUT11), .ZN(new_n518_));
  XOR2_X1   g317(.A(G71gat), .B(G78gat), .Z(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n518_), .A2(new_n519_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n507_), .A2(new_n515_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n492_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n492_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT67), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n515_), .B(KEYINPUT66), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n507_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n522_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT12), .A3(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n525_), .B2(KEYINPUT12), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n526_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT70), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G120gat), .B(G148gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G176gat), .B(G204gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n535_), .A2(new_n543_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT13), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n537_), .A2(new_n548_), .A3(new_n545_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n531_), .A2(new_n466_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n507_), .A2(new_n515_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n465_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT73), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI22_X1  g363(.A1(new_n558_), .A2(new_n559_), .B1(KEYINPUT35), .B2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n557_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT74), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(KEYINPUT35), .ZN(new_n569_));
  OR3_X1    g368(.A1(new_n566_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n566_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(KEYINPUT36), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n570_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT75), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT75), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n570_), .A2(new_n571_), .A3(new_n578_), .A4(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT37), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n570_), .A2(new_n571_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n574_), .B(KEYINPUT36), .Z(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n570_), .A2(new_n571_), .A3(KEYINPUT76), .ZN(new_n586_));
  INV_X1    g385(.A(new_n583_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT76), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n586_), .A2(new_n589_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n585_), .B1(new_n590_), .B2(KEYINPUT37), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n473_), .B(new_n522_), .Z(new_n592_));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  OR3_X1    g398(.A1(new_n594_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(KEYINPUT17), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n594_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n591_), .A2(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n490_), .A2(new_n556_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n428_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  AOI21_X1  g407(.A(G1gat), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n607_), .A2(new_n608_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n442_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n451_), .A2(new_n452_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n429_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT100), .B1(new_n615_), .B2(new_n443_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n613_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n589_), .A2(new_n586_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n580_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n489_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n603_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n556_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT102), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(new_n606_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n612_), .B1(new_n626_), .B2(new_n468_), .ZN(G1324gat));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628_));
  INV_X1    g427(.A(new_n459_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(KEYINPUT103), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G8gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT103), .B1(new_n624_), .B2(new_n629_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT104), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(G8gat), .A4(new_n630_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n633_), .A2(new_n636_), .A3(KEYINPUT39), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n605_), .A2(new_n469_), .A3(new_n629_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(new_n633_), .B2(KEYINPUT39), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n628_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n633_), .A2(new_n636_), .A3(KEYINPUT39), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n641_), .A2(KEYINPUT40), .A3(new_n642_), .A4(new_n638_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n625_), .B2(new_n248_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT41), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n605_), .A2(new_n645_), .A3(new_n248_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1326gat));
  INV_X1    g448(.A(G22gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n421_), .B(KEYINPUT105), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n625_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT42), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n605_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1327gat));
  AOI21_X1  g454(.A(KEYINPUT107), .B1(new_n590_), .B2(new_n603_), .ZN(new_n656_));
  AND4_X1   g455(.A1(KEYINPUT107), .A2(new_n618_), .A3(new_n580_), .A4(new_n603_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n555_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n553_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n490_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G29gat), .B1(new_n663_), .B2(new_n606_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n659_), .A2(new_n621_), .A3(new_n553_), .A4(new_n603_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT106), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n617_), .A2(new_n667_), .A3(new_n591_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n619_), .A2(new_n581_), .B1(new_n580_), .B2(new_n584_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT43), .B1(new_n461_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT44), .B1(new_n666_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n666_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n606_), .A2(G29gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n664_), .B1(new_n675_), .B2(new_n676_), .ZN(G1328gat));
  OR2_X1    g476(.A1(new_n629_), .A2(KEYINPUT108), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n629_), .A2(KEYINPUT108), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n662_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n662_), .A2(KEYINPUT45), .A3(new_n682_), .ZN(new_n686_));
  OAI22_X1  g485(.A1(new_n685_), .A2(new_n686_), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n673_), .A2(new_n629_), .A3(new_n674_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(G36gat), .B2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1329gat));
  NOR2_X1   g490(.A1(new_n246_), .A2(new_n242_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n675_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G43gat), .B1(new_n663_), .B2(new_n248_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT47), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n693_), .A2(new_n698_), .A3(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1330gat));
  AOI21_X1  g499(.A(G50gat), .B1(new_n663_), .B2(new_n651_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n429_), .A2(G50gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n675_), .B2(new_n702_), .ZN(G1331gat));
  NOR2_X1   g502(.A1(new_n603_), .A2(new_n621_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n617_), .A2(new_n619_), .A3(new_n660_), .A4(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT112), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(G57gat), .A3(new_n606_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT113), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT113), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n604_), .A2(new_n660_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT110), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n617_), .A2(new_n715_), .A3(new_n489_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT111), .B1(new_n461_), .B2(new_n621_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n714_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n606_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n711_), .A2(new_n712_), .A3(new_n721_), .ZN(G1332gat));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n723_), .A3(new_n680_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n709_), .A2(new_n680_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(G64gat), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT48), .B(new_n723_), .C1(new_n709_), .C2(new_n680_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n720_), .A2(new_n730_), .A3(new_n248_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT49), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n709_), .A2(new_n248_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G71gat), .ZN(new_n734_));
  AOI211_X1 g533(.A(KEYINPUT49), .B(new_n730_), .C1(new_n709_), .C2(new_n248_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n720_), .A2(new_n737_), .A3(new_n651_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n707_), .A2(new_n651_), .A3(new_n708_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(new_n740_), .A3(G78gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n739_), .B2(G78gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(G1335gat));
  OAI22_X1  g544(.A1(new_n657_), .A2(new_n656_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n715_), .B1(new_n617_), .B2(new_n489_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n461_), .A2(KEYINPUT111), .A3(new_n621_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT115), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n718_), .A2(new_n752_), .A3(new_n747_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n512_), .A3(new_n606_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n489_), .B(new_n603_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n428_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n759_), .ZN(G1336gat));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n513_), .A3(new_n629_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n680_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G92gat), .B1(new_n758_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1337gat));
  INV_X1    g563(.A(new_n508_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n246_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n248_), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n769_), .B(new_n756_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n770_));
  INV_X1    g569(.A(G99gat), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n768_), .B2(new_n772_), .ZN(new_n773_));
  XOR2_X1   g572(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n768_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n752_), .B1(new_n718_), .B2(new_n747_), .ZN(new_n779_));
  AOI211_X1 g578(.A(KEYINPUT115), .B(new_n746_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n766_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n757_), .A2(new_n248_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n774_), .B1(new_n782_), .B2(G99gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT117), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n773_), .B1(new_n778_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT118), .B(new_n773_), .C1(new_n778_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n754_), .A2(new_n509_), .A3(new_n429_), .ZN(new_n790_));
  AOI211_X1 g589(.A(KEYINPUT52), .B(new_n509_), .C1(new_n757_), .C2(new_n429_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n757_), .A2(new_n429_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(G106gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n475_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n479_), .A2(new_n477_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n487_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n487_), .B2(new_n482_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n550_), .A2(new_n552_), .A3(new_n801_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n534_), .A2(new_n524_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n492_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n529_), .A2(new_n807_), .A3(new_n534_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n803_), .A2(KEYINPUT119), .A3(new_n492_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n806_), .A2(new_n808_), .A3(new_n809_), .A4(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT120), .B1(new_n811_), .B2(new_n543_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(KEYINPUT56), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n547_), .A2(new_n489_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n812_), .B2(KEYINPUT56), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n802_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n619_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n820_));
  OR2_X1    g619(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n811_), .A2(new_n543_), .A3(new_n820_), .A4(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n547_), .A2(new_n800_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n811_), .A2(new_n543_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n822_), .B(new_n823_), .C1(new_n824_), .C2(new_n820_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n669_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n825_), .A2(new_n826_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n819_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n817_), .A2(new_n818_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n603_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n604_), .A2(new_n556_), .A3(new_n489_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT54), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n428_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(G113gat), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n629_), .A2(new_n429_), .A3(new_n246_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n621_), .A4(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(KEYINPUT59), .A3(new_n837_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n831_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n817_), .A2(new_n818_), .B1(new_n828_), .B2(new_n827_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n622_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n834_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n606_), .B(new_n837_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n489_), .B1(new_n839_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n838_), .B1(new_n847_), .B2(new_n836_), .ZN(G1340gat));
  XOR2_X1   g647(.A(KEYINPUT122), .B(G120gat), .Z(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n556_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(KEYINPUT60), .B2(new_n849_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n844_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n556_), .B1(new_n839_), .B2(new_n846_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n849_), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n835_), .A2(new_n855_), .A3(new_n622_), .A4(new_n837_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n603_), .B1(new_n839_), .B2(new_n846_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n855_), .ZN(G1342gat));
  NAND2_X1  g657(.A1(new_n839_), .A2(new_n846_), .ZN(new_n859_));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n669_), .A2(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT123), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n835_), .A2(new_n590_), .A3(new_n837_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n859_), .A2(new_n862_), .B1(new_n863_), .B2(new_n860_), .ZN(G1343gat));
  NOR3_X1   g663(.A1(new_n680_), .A2(new_n421_), .A3(new_n248_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n835_), .A2(new_n621_), .A3(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT124), .B(G141gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n835_), .A2(new_n660_), .A3(new_n865_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g669(.A1(new_n835_), .A2(new_n622_), .A3(new_n865_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  NAND2_X1  g672(.A1(new_n835_), .A2(new_n865_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G162gat), .B1(new_n874_), .B2(new_n669_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n619_), .A2(G162gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n874_), .B2(new_n876_), .ZN(G1347gat));
  NAND2_X1  g676(.A1(new_n832_), .A2(new_n834_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n680_), .A2(new_n428_), .A3(new_n248_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n651_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n621_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(G169gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(G169gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n878_), .A2(new_n880_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n621_), .A2(new_n221_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT125), .ZN(new_n887_));
  OAI22_X1  g686(.A1(new_n883_), .A2(new_n884_), .B1(new_n885_), .B2(new_n887_), .ZN(G1348gat));
  INV_X1    g687(.A(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n660_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n429_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n879_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(G176gat), .A3(new_n660_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n890_), .A2(new_n222_), .B1(new_n891_), .B2(new_n894_), .ZN(G1349gat));
  NOR3_X1   g694(.A1(new_n885_), .A2(new_n203_), .A3(new_n603_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n891_), .A2(new_n622_), .A3(new_n892_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n225_), .B2(new_n897_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n885_), .B2(new_n669_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n590_), .A2(new_n204_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n885_), .B2(new_n900_), .ZN(G1351gat));
  NOR4_X1   g700(.A1(new_n762_), .A2(new_n606_), .A3(new_n421_), .A4(new_n248_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n878_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n489_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n285_), .ZN(G1352gat));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n556_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(KEYINPUT126), .B2(new_n286_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT126), .B(G204gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(new_n908_), .ZN(G1353gat));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n622_), .B1(new_n910_), .B2(new_n294_), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT127), .Z(new_n912_));
  NOR2_X1   g711(.A1(new_n903_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1354gat));
  OAI21_X1  g714(.A(G218gat), .B1(new_n903_), .B2(new_n669_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n590_), .A2(new_n292_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n903_), .B2(new_n917_), .ZN(G1355gat));
endmodule


