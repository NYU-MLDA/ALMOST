//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_;
  INV_X1    g000(.A(KEYINPUT106), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT79), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT22), .B(G169gat), .Z(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT95), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT81), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT82), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(new_n213_), .B2(KEYINPUT23), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n220_));
  OAI22_X1  g019(.A1(new_n217_), .A2(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n213_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT23), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n214_), .B2(KEYINPUT23), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  AOI211_X1 g028(.A(new_n225_), .B(new_n227_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n212_), .A2(new_n221_), .B1(new_n224_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G197gat), .B(G204gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT21), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n233_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n237_), .A3(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT20), .B1(new_n231_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n214_), .A2(new_n215_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n219_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n225_), .B1(new_n244_), .B2(new_n216_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n246_));
  INV_X1    g045(.A(G183gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT25), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n247_), .A2(KEYINPUT25), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n228_), .B(new_n248_), .C1(new_n249_), .C2(new_n246_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n208_), .B2(new_n226_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT80), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT80), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n250_), .B(new_n253_), .C1(new_n208_), .C2(new_n226_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n245_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n224_), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n208_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT83), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT22), .B1(new_n258_), .B2(G169gat), .ZN(new_n259_));
  INV_X1    g058(.A(G169gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT84), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT22), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(KEYINPUT83), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n211_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n256_), .B(new_n257_), .C1(new_n262_), .C2(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n255_), .A2(new_n240_), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n206_), .B1(new_n241_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n269_), .B1(new_n231_), .B2(new_n240_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n255_), .A2(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n239_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n272_), .A3(new_n205_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G8gat), .B(G36gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n268_), .A2(new_n279_), .A3(new_n273_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(KEYINPUT97), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n274_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT97), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(new_n279_), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n241_), .A2(new_n267_), .A3(new_n206_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n205_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n280_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT27), .A3(new_n282_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT3), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT2), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n301_), .B1(KEYINPUT1), .B2(new_n303_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(KEYINPUT1), .B2(new_n303_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n296_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n307_), .A2(new_n298_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n300_), .A2(new_n304_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310_));
  XOR2_X1   g109(.A(G22gat), .B(G50gat), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n295_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n294_), .A3(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G228gat), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT89), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n300_), .A2(new_n304_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n306_), .A2(new_n308_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n324_), .B1(new_n327_), .B2(KEYINPUT29), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n309_), .A2(new_n323_), .A3(new_n310_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n239_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(KEYINPUT29), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT89), .B1(new_n236_), .B2(new_n238_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n320_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n330_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n319_), .B(new_n336_), .C1(new_n337_), .C2(KEYINPUT92), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n330_), .A2(new_n334_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n335_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(KEYINPUT92), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n327_), .A2(KEYINPUT90), .A3(KEYINPUT29), .ZN(new_n343_));
  INV_X1    g142(.A(new_n324_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n240_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n321_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n340_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n319_), .B1(new_n336_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT91), .ZN(new_n350_));
  OAI22_X1  g149(.A1(new_n338_), .A2(new_n342_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n350_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT93), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n349_), .A2(new_n350_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT92), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n341_), .A2(new_n357_), .A3(new_n319_), .A4(new_n336_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT93), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n355_), .A2(new_n352_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n293_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT100), .ZN(new_n364_));
  INV_X1    g163(.A(G1gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n367_));
  INV_X1    g166(.A(G29gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n366_), .B(new_n369_), .Z(new_n370_));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n372_), .A2(KEYINPUT86), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(KEYINPUT86), .ZN(new_n374_));
  XOR2_X1   g173(.A(G113gat), .B(G120gat), .Z(new_n375_));
  OR3_X1    g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n309_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n371_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n377_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n327_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n309_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT4), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT98), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n380_), .A2(new_n384_), .A3(KEYINPUT98), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n382_), .A2(new_n383_), .A3(new_n371_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n370_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n366_), .B(new_n369_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n387_), .A2(new_n393_), .A3(new_n390_), .A4(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G71gat), .B(G99gat), .ZN(new_n396_));
  INV_X1    g195(.A(G43gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(G15gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n398_), .B(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n255_), .A2(KEYINPUT30), .A3(new_n266_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT30), .B1(new_n255_), .B2(new_n266_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT85), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n403_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n402_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n402_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n381_), .B(KEYINPUT31), .Z(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n412_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n410_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n362_), .A2(new_n395_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n382_), .A2(new_n383_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n370_), .B1(new_n420_), .B2(new_n371_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n378_), .A2(new_n379_), .B1(G225gat), .B2(G233gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n384_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n394_), .A2(KEYINPUT33), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n389_), .A2(new_n390_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n393_), .A4(new_n387_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n282_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n279_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n285_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n274_), .A2(KEYINPUT97), .A3(new_n280_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n428_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n279_), .A2(KEYINPUT32), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT101), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n284_), .A2(KEYINPUT102), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n268_), .A2(new_n435_), .A3(new_n273_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT102), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT32), .B(new_n279_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n395_), .A2(new_n436_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n433_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n395_), .B1(new_n354_), .B2(new_n360_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n361_), .A2(new_n442_), .B1(new_n293_), .B2(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n414_), .A2(KEYINPUT87), .A3(new_n417_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT87), .B1(new_n414_), .B2(new_n417_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT104), .B1(new_n444_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n442_), .A2(new_n361_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n354_), .A2(new_n360_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n395_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n288_), .A4(new_n292_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT104), .ZN(new_n454_));
  INV_X1    g253(.A(new_n447_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n419_), .B1(new_n448_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G8gat), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT76), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(KEYINPUT76), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n365_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n459_), .A2(new_n464_), .A3(new_n462_), .A4(new_n460_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n468_), .B(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G229gat), .A2(G233gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n471_), .B(KEYINPUT15), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n467_), .A3(new_n466_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n472_), .A2(new_n474_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G113gat), .B(G141gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G169gat), .B(G197gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  XOR2_X1   g280(.A(new_n478_), .B(new_n481_), .Z(new_n482_));
  NOR2_X1   g281(.A1(new_n457_), .A2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(G71gat), .A2(G78gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G71gat), .A2(G78gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G57gat), .B(G64gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(KEYINPUT11), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n487_), .B2(KEYINPUT11), .ZN(new_n490_));
  INV_X1    g289(.A(G64gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G57gat), .ZN(new_n492_));
  INV_X1    g291(.A(G57gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G64gat), .ZN(new_n494_));
  AND4_X1   g293(.A1(new_n489_), .A2(new_n492_), .A3(new_n494_), .A4(KEYINPUT11), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n488_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n494_), .A3(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT68), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n492_), .A2(new_n494_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT11), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n492_), .A2(new_n494_), .A3(new_n489_), .A4(KEYINPUT11), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n498_), .A2(new_n501_), .A3(new_n486_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n496_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n507_));
  INV_X1    g306(.A(G99gat), .ZN(new_n508_));
  INV_X1    g307(.A(G106gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT7), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT6), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT7), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n507_), .A2(new_n517_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n511_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT8), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n519_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT9), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G85gat), .ZN(new_n529_));
  INV_X1    g328(.A(G92gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT65), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT65), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(G92gat), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n529_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n520_), .A2(new_n521_), .A3(new_n528_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT66), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G85gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT9), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n532_), .A2(G92gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n530_), .A2(KEYINPUT65), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT66), .ZN(new_n542_));
  INV_X1    g341(.A(new_n521_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(KEYINPUT9), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n536_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT10), .B(G99gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n516_), .B1(new_n549_), .B2(G106gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n527_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n536_), .B2(new_n546_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(new_n548_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n506_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n524_), .A2(new_n526_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n505_), .B1(new_n557_), .B2(new_n504_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT64), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n557_), .B2(new_n504_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT70), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n557_), .A2(new_n504_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT66), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n542_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n551_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n525_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n519_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n569_), .B(new_n504_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n561_), .B1(new_n566_), .B2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n556_), .A2(KEYINPUT70), .A3(new_n558_), .A4(new_n562_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n565_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT5), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n565_), .A2(new_n574_), .A3(new_n575_), .A4(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT71), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT13), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n581_), .B(new_n583_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n583_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n589_));
  OAI21_X1  g388(.A(new_n586_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT72), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(KEYINPUT74), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n599_));
  OAI22_X1  g398(.A1(new_n596_), .A2(new_n599_), .B1(KEYINPUT35), .B2(new_n593_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n471_), .B2(new_n557_), .ZN(new_n601_));
  OAI211_X1 g400(.A(KEYINPUT73), .B(new_n475_), .C1(new_n553_), .C2(new_n555_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n548_), .A2(new_n554_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n569_), .A2(KEYINPUT69), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT73), .B1(new_n606_), .B2(new_n475_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n598_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n475_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT73), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n598_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n602_), .A4(new_n601_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT36), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT75), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n608_), .A2(new_n613_), .A3(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n616_), .A2(KEYINPUT36), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n608_), .B2(new_n613_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT37), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n608_), .A2(new_n613_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n620_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT37), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n608_), .A2(new_n613_), .A3(new_n618_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n468_), .B(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n504_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n504_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT17), .ZN(new_n635_));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT16), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G183gat), .B(G211gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  OAI22_X1  g438(.A1(new_n633_), .A2(new_n634_), .B1(new_n635_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n634_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n639_), .B(new_n635_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n632_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT77), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n640_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n629_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n591_), .A2(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n483_), .A2(new_n365_), .A3(new_n395_), .A4(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(KEYINPUT38), .A3(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n619_), .A2(new_n622_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n482_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n590_), .A2(new_n656_), .A3(new_n648_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n457_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n395_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G1gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n654_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT38), .B1(new_n652_), .B2(new_n653_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n202_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n662_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n664_), .A2(KEYINPUT106), .A3(new_n660_), .A4(new_n654_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1324gat));
  XNOR2_X1  g465(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n669_));
  INV_X1    g468(.A(new_n419_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n454_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT104), .B(new_n447_), .C1(new_n449_), .C2(new_n452_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n293_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n655_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n657_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G8gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n669_), .B1(new_n678_), .B2(KEYINPUT39), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n677_), .A2(KEYINPUT108), .A3(new_n680_), .A4(G8gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT107), .B(new_n680_), .C1(new_n677_), .C2(G8gat), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n678_), .B2(KEYINPUT39), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n682_), .A2(new_n683_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n483_), .A2(new_n650_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n687_), .A2(G8gat), .A3(new_n293_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n668_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n688_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n685_), .A2(new_n683_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n690_), .B(new_n667_), .C1(new_n691_), .C2(new_n682_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(G1325gat));
  INV_X1    g492(.A(new_n687_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n400_), .A3(new_n447_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n658_), .A2(new_n447_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n696_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT41), .B1(new_n696_), .B2(G15gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n695_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT110), .Z(G1326gat));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n450_), .B(KEYINPUT111), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n658_), .B2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT42), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n694_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1327gat));
  NOR3_X1   g506(.A1(new_n591_), .A2(new_n648_), .A3(new_n675_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n483_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n395_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n457_), .B2(new_n629_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n623_), .A2(new_n628_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n673_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n590_), .A2(new_n656_), .A3(new_n647_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT44), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n719_), .B(new_n716_), .C1(new_n711_), .C2(new_n714_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n451_), .A2(new_n368_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n710_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(KEYINPUT46), .ZN(new_n725_));
  INV_X1    g524(.A(G36gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n721_), .B2(new_n674_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n709_), .A2(new_n726_), .A3(new_n674_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n725_), .B1(new_n727_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n728_), .B(KEYINPUT45), .ZN(new_n732_));
  INV_X1    g531(.A(new_n725_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n718_), .A2(new_n720_), .A3(new_n293_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n732_), .B(new_n733_), .C1(new_n726_), .C2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n735_), .ZN(G1329gat));
  AOI21_X1  g535(.A(G43gat), .B1(new_n709_), .B2(new_n447_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n418_), .A2(new_n397_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n721_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1330gat));
  INV_X1    g540(.A(G50gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n709_), .A2(new_n742_), .A3(new_n703_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n721_), .A2(KEYINPUT113), .A3(new_n450_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G50gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT113), .B1(new_n721_), .B2(new_n450_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n745_), .B2(new_n746_), .ZN(G1331gat));
  NOR4_X1   g546(.A1(new_n457_), .A2(new_n656_), .A3(new_n590_), .A4(new_n649_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n493_), .A3(new_n395_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n590_), .A2(new_n656_), .A3(new_n647_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n673_), .A2(new_n675_), .A3(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G57gat), .B1(new_n751_), .B2(new_n451_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1332gat));
  NAND3_X1  g552(.A1(new_n748_), .A2(new_n491_), .A3(new_n674_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G64gat), .B1(new_n751_), .B2(new_n293_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n755_), .A2(new_n757_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT115), .Z(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n751_), .B2(new_n455_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  INV_X1    g562(.A(G71gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n748_), .A2(new_n764_), .A3(new_n447_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1334gat));
  OAI21_X1  g565(.A(G78gat), .B1(new_n751_), .B2(new_n702_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT50), .ZN(new_n768_));
  INV_X1    g567(.A(G78gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n748_), .A2(new_n769_), .A3(new_n703_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1335gat));
  NAND3_X1  g570(.A1(new_n591_), .A2(new_n482_), .A3(new_n647_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT116), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n451_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n590_), .A2(new_n648_), .A3(new_n675_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n673_), .A2(new_n482_), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n537_), .A3(new_n395_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(G1336gat));
  AOI21_X1  g579(.A(G92gat), .B1(new_n778_), .B2(new_n674_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n293_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n774_), .B2(new_n782_), .ZN(G1337gat));
  AOI21_X1  g582(.A(new_n508_), .B1(new_n774_), .B2(new_n447_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n418_), .A2(new_n549_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n778_), .B2(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g586(.A1(new_n778_), .A2(new_n509_), .A3(new_n450_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n774_), .A2(new_n450_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G106gat), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT52), .B(new_n509_), .C1(new_n774_), .C2(new_n450_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n788_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n481_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n473_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n476_), .A2(new_n800_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n478_), .A2(new_n481_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n583_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n565_), .A2(new_n804_), .A3(new_n575_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n496_), .A2(new_n503_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT12), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n567_), .A2(new_n568_), .ZN(new_n809_));
  OAI22_X1  g608(.A1(new_n809_), .A2(new_n550_), .B1(new_n571_), .B2(new_n570_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT12), .B1(new_n810_), .B2(new_n806_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n572_), .A2(new_n560_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n808_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n556_), .A2(new_n572_), .A3(new_n558_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n813_), .A2(KEYINPUT55), .B1(new_n814_), .B2(new_n561_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n805_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n580_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n580_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n803_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n713_), .B1(new_n821_), .B2(KEYINPUT58), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(KEYINPUT58), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT117), .B(new_n713_), .C1(new_n821_), .C2(KEYINPUT58), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n816_), .B2(new_n580_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n818_), .B(new_n582_), .C1(new_n805_), .C2(new_n815_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n656_), .B(new_n583_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n587_), .A2(new_n802_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT57), .B1(new_n832_), .B2(new_n675_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n834_), .B(new_n655_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n648_), .B1(new_n827_), .B2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n590_), .A2(new_n629_), .A3(new_n482_), .A4(new_n648_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n798_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n656_), .A2(new_n583_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n831_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n675_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n834_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n832_), .A2(KEYINPUT57), .A3(new_n675_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n826_), .A2(new_n825_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n803_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT117), .B1(new_n852_), .B2(new_n713_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n846_), .B(new_n847_), .C1(new_n848_), .C2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n647_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n840_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(KEYINPUT118), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n841_), .A2(new_n857_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n362_), .A2(new_n451_), .A3(new_n418_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT59), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n862_), .B(new_n859_), .C1(new_n837_), .C2(new_n840_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n656_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G113gat), .ZN(new_n866_));
  OR3_X1    g665(.A1(new_n860_), .A2(G113gat), .A3(new_n482_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(new_n860_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n590_), .A2(KEYINPUT60), .ZN(new_n870_));
  MUX2_X1   g669(.A(new_n870_), .B(KEYINPUT60), .S(G120gat), .Z(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n861_), .A2(new_n591_), .A3(new_n863_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT119), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G120gat), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(KEYINPUT119), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n872_), .B1(new_n875_), .B2(new_n876_), .ZN(G1341gat));
  NAND2_X1  g676(.A1(new_n864_), .A2(new_n648_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G127gat), .ZN(new_n879_));
  OR3_X1    g678(.A1(new_n860_), .A2(G127gat), .A3(new_n647_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1342gat));
  AOI21_X1  g680(.A(G134gat), .B1(new_n869_), .B2(new_n655_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT120), .B(G134gat), .Z(new_n883_));
  NOR2_X1   g682(.A1(new_n629_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n864_), .B2(new_n884_), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n361_), .A2(new_n451_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n455_), .A2(new_n886_), .A3(new_n293_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT118), .B1(new_n855_), .B2(new_n856_), .ZN(new_n889_));
  AOI211_X1 g688(.A(new_n798_), .B(new_n840_), .C1(new_n854_), .C2(new_n647_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT121), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n858_), .A2(new_n893_), .A3(new_n888_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n656_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n591_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n895_), .B2(new_n648_), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT122), .B(new_n647_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n901_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n893_), .B1(new_n858_), .B2(new_n888_), .ZN(new_n906_));
  AOI211_X1 g705(.A(KEYINPUT121), .B(new_n887_), .C1(new_n841_), .C2(new_n857_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n648_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT122), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n895_), .A2(new_n902_), .A3(new_n648_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n910_), .A3(new_n900_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n905_), .A2(new_n911_), .ZN(G1346gat));
  INV_X1    g711(.A(G162gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n895_), .A2(new_n913_), .A3(new_n655_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n629_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n913_), .ZN(G1347gat));
  AOI21_X1  g715(.A(new_n703_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n455_), .A2(new_n395_), .A3(new_n293_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n656_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n921_), .A2(new_n922_), .A3(G169gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n921_), .B2(G169gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n656_), .A2(new_n210_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT123), .ZN(new_n927_));
  OAI22_X1  g726(.A1(new_n924_), .A2(new_n925_), .B1(new_n919_), .B2(new_n927_), .ZN(G1348gat));
  AOI21_X1  g727(.A(G176gat), .B1(new_n920_), .B2(new_n591_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n590_), .A2(new_n211_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n858_), .A2(new_n361_), .A3(new_n918_), .A4(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n932_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n929_), .B1(new_n933_), .B2(new_n934_), .ZN(G1349gat));
  NAND4_X1  g734(.A1(new_n858_), .A2(new_n361_), .A3(new_n648_), .A4(new_n918_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n918_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n937_), .A2(new_n229_), .A3(new_n647_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n936_), .A2(new_n247_), .B1(new_n917_), .B2(new_n938_), .ZN(G1350gat));
  OAI21_X1  g738(.A(G190gat), .B1(new_n919_), .B2(new_n629_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n655_), .A2(new_n228_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n919_), .B2(new_n941_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT125), .ZN(G1351gat));
  NOR4_X1   g742(.A1(new_n447_), .A2(new_n293_), .A3(new_n361_), .A4(new_n395_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n858_), .A2(new_n944_), .ZN(new_n945_));
  OR2_X1    g744(.A1(new_n945_), .A2(KEYINPUT126), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(KEYINPUT126), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(G197gat), .B1(new_n948_), .B2(new_n656_), .ZN(new_n949_));
  INV_X1    g748(.A(G197gat), .ZN(new_n950_));
  AOI211_X1 g749(.A(new_n950_), .B(new_n482_), .C1(new_n946_), .C2(new_n947_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n949_), .A2(new_n951_), .ZN(G1352gat));
  NAND2_X1  g751(.A1(new_n948_), .A2(new_n591_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(G204gat), .ZN(new_n954_));
  INV_X1    g753(.A(G204gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n948_), .A2(new_n955_), .A3(new_n591_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n956_), .ZN(G1353gat));
  NOR2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(KEYINPUT127), .ZN(new_n959_));
  NAND2_X1  g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n648_), .A2(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n959_), .B1(new_n948_), .B2(new_n962_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n959_), .ZN(new_n964_));
  AOI211_X1 g763(.A(new_n964_), .B(new_n961_), .C1(new_n946_), .C2(new_n947_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n963_), .A2(new_n965_), .ZN(G1354gat));
  INV_X1    g765(.A(G218gat), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n948_), .A2(new_n967_), .A3(new_n655_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n629_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n967_), .ZN(G1355gat));
endmodule


