//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT85), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n205_), .A2(KEYINPUT1), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(KEYINPUT1), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT86), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(KEYINPUT86), .A3(KEYINPUT1), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n206_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT84), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT84), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n204_), .A2(new_n219_), .A3(new_n205_), .ZN(new_n220_));
  INV_X1    g019(.A(G155gat), .ZN(new_n221_));
  INV_X1    g020(.A(G162gat), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT85), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT85), .B1(new_n221_), .B2(new_n222_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n205_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT87), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n213_), .A2(new_n215_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n217_), .A2(KEYINPUT3), .ZN(new_n230_));
  OR3_X1    g029(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n220_), .A2(new_n226_), .A3(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n218_), .A2(new_n233_), .A3(KEYINPUT88), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT88), .B1(new_n218_), .B2(new_n233_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G22gat), .B(G50gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT28), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n202_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n240_), .A3(KEYINPUT89), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G211gat), .B(G218gat), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT92), .B1(new_n247_), .B2(G197gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(KEYINPUT21), .A3(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G197gat), .B(G204gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n246_), .A2(KEYINPUT21), .ZN(new_n252_));
  XOR2_X1   g051(.A(G197gat), .B(G204gat), .Z(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(KEYINPUT21), .A3(new_n246_), .A4(new_n248_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G228gat), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT90), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(KEYINPUT90), .ZN(new_n259_));
  AND2_X1   g058(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n258_), .B(new_n259_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n256_), .B(new_n262_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G78gat), .B(G106gat), .Z(new_n264_));
  INV_X1    g063(.A(new_n262_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(KEYINPUT93), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT93), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n251_), .A2(new_n254_), .A3(new_n267_), .A4(new_n252_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n237_), .B1(new_n218_), .B2(new_n233_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n265_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n263_), .A2(new_n264_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n264_), .B1(new_n263_), .B2(new_n271_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n243_), .B(new_n245_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n241_), .A2(new_n242_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n263_), .A2(new_n271_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n264_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n275_), .B1(new_n278_), .B2(KEYINPUT94), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n263_), .A2(new_n264_), .A3(new_n271_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT94), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(new_n273_), .B2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n274_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT23), .ZN(new_n287_));
  INV_X1    g086(.A(G169gat), .ZN(new_n288_));
  INV_X1    g087(.A(G176gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT24), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n287_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT80), .B(G183gat), .Z(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(KEYINPUT25), .ZN(new_n297_));
  NOR2_X1   g096(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT81), .B(G190gat), .Z(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(KEYINPUT26), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n294_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n287_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT22), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT82), .B1(new_n303_), .B2(G169gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n289_), .B(new_n304_), .C1(new_n305_), .C2(KEYINPUT82), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n292_), .A3(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n301_), .A2(new_n255_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n287_), .B1(G183gat), .B2(G190gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n289_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n292_), .B(KEYINPUT97), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT96), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n287_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT25), .B(G183gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT26), .B(G190gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n294_), .A2(KEYINPUT96), .A3(new_n317_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n312_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(KEYINPUT20), .B(new_n308_), .C1(new_n321_), .C2(new_n255_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT95), .Z(new_n324_));
  XOR2_X1   g123(.A(new_n324_), .B(KEYINPUT19), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT18), .B(G64gat), .ZN(new_n328_));
  INV_X1    g127(.A(G92gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n321_), .A2(new_n255_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT20), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n301_), .A2(new_n307_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n256_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n325_), .A3(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n327_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n327_), .B2(new_n337_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n285_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n327_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n322_), .A2(new_n326_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n312_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n269_), .B(new_n343_), .C1(new_n314_), .C2(new_n318_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n325_), .B1(new_n344_), .B2(new_n336_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(KEYINPUT27), .B(new_n341_), .C1(new_n346_), .C2(new_n332_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n340_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n284_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n335_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n352_), .B(KEYINPUT30), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n351_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G71gat), .B(G99gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n354_), .B(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G127gat), .B(G134gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G113gat), .ZN(new_n359_));
  INV_X1    g158(.A(G120gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G15gat), .B(G43gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT31), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n361_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n357_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT0), .B(G57gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G85gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(G1gat), .B(G29gat), .Z(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n218_), .A2(new_n233_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n218_), .A2(new_n233_), .A3(KEYINPUT88), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n361_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n359_), .B(G120gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(new_n371_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT4), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n370_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n361_), .A2(new_n233_), .A3(new_n218_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n370_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n369_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n380_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n373_), .A2(new_n374_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT4), .B1(new_n389_), .B2(new_n376_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n384_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n370_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n369_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n387_), .A2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n349_), .A2(new_n365_), .A3(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n387_), .A2(new_n395_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n283_), .A2(new_n348_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT100), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n283_), .A2(new_n398_), .A3(new_n348_), .A4(KEYINPUT100), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n327_), .A2(new_n337_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n346_), .A2(new_n403_), .ZN(new_n406_));
  AOI211_X1 g205(.A(new_n405_), .B(new_n406_), .C1(new_n387_), .C2(new_n395_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT98), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n395_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n395_), .B2(new_n408_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n370_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT99), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n394_), .B1(new_n392_), .B2(new_n385_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n416_), .B(new_n370_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n338_), .A2(new_n339_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n407_), .B1(new_n412_), .B2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n401_), .B(new_n402_), .C1(new_n421_), .C2(new_n283_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n397_), .B1(new_n422_), .B2(new_n365_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT16), .B(G183gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G211gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G127gat), .B(G155gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT66), .B1(new_n427_), .B2(KEYINPUT17), .ZN(new_n428_));
  OR2_X1    g227(.A1(G71gat), .A2(G78gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G71gat), .A2(G78gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(G57gat), .A2(G64gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G57gat), .A2(G64gat), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n433_), .A2(new_n434_), .A3(KEYINPUT11), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT11), .ZN(new_n436_));
  INV_X1    g235(.A(G57gat), .ZN(new_n437_));
  INV_X1    g236(.A(G64gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G57gat), .A2(G64gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n436_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n432_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT11), .B1(new_n433_), .B2(new_n434_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n431_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G15gat), .B(G22gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G1gat), .A2(G8gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT14), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G1gat), .ZN(new_n450_));
  INV_X1    g249(.A(G8gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n447_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n446_), .A2(new_n447_), .A3(new_n452_), .A4(new_n448_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n445_), .B(new_n456_), .Z(new_n457_));
  XNOR2_X1  g256(.A(new_n428_), .B(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G231gat), .A2(G233gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n459_), .B(KEYINPUT78), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n458_), .B(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n427_), .A2(KEYINPUT17), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n423_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n466_));
  INV_X1    g265(.A(G99gat), .ZN(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n469_), .A2(new_n472_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n329_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT8), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT8), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n472_), .A2(new_n473_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(KEYINPUT9), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT9), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT65), .B1(new_n478_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n486_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n467_), .A2(KEYINPUT10), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT10), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G99gat), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n491_), .A2(new_n493_), .A3(KEYINPUT64), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT64), .B1(new_n491_), .B2(new_n493_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n468_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n482_), .A2(new_n484_), .B1(new_n490_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT66), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n442_), .A2(new_n498_), .A3(new_n444_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n439_), .A2(new_n436_), .A3(new_n440_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n431_), .B1(new_n443_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n439_), .A2(new_n440_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n502_), .A2(KEYINPUT11), .B1(new_n429_), .B2(new_n430_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT66), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT67), .B1(new_n497_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n497_), .A2(new_n505_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n497_), .B2(new_n505_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n445_), .A2(KEYINPUT12), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n514_), .B1(new_n497_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n497_), .A2(new_n505_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n475_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n483_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT64), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n492_), .A2(G99gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n467_), .A2(KEYINPUT10), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n491_), .A2(new_n493_), .A3(KEYINPUT64), .ZN(new_n524_));
  AOI21_X1  g323(.A(G106gat), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n473_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n488_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n478_), .A2(new_n488_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT65), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n528_), .B(new_n485_), .C1(new_n529_), .C2(new_n532_), .ZN(new_n533_));
  OAI22_X1  g332(.A1(new_n518_), .A2(new_n519_), .B1(new_n525_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n512_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT68), .A3(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n513_), .A2(new_n516_), .A3(new_n517_), .A4(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n511_), .B1(new_n510_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n247_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT5), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(new_n289_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT69), .Z(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n511_), .B(new_n542_), .C1(new_n510_), .C2(new_n537_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n538_), .A2(KEYINPUT70), .A3(new_n543_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT13), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G43gat), .B(G50gat), .ZN(new_n553_));
  INV_X1    g352(.A(G29gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT71), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT71), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G29gat), .ZN(new_n557_));
  INV_X1    g356(.A(G36gat), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n555_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n553_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n556_), .A2(G29gat), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n554_), .A2(KEYINPUT71), .ZN(new_n563_));
  OAI21_X1  g362(.A(G36gat), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G43gat), .B(G50gat), .Z(new_n565_));
  NAND3_X1  g364(.A1(new_n555_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n456_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n561_), .A2(new_n567_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n552_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n559_), .A2(new_n560_), .A3(new_n553_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n565_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n561_), .A2(new_n567_), .A3(KEYINPUT15), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n572_), .B1(new_n578_), .B2(new_n456_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n571_), .B1(new_n579_), .B2(new_n552_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(new_n288_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G197gat), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n580_), .A2(KEYINPUT79), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT79), .B1(new_n580_), .B2(new_n583_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n580_), .A2(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n551_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n465_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT35), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n497_), .A2(new_n567_), .A3(new_n561_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n561_), .A2(KEYINPUT15), .A3(new_n567_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT15), .B1(new_n561_), .B2(new_n567_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n534_), .B(new_n599_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n599_), .B1(new_n578_), .B2(new_n534_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n597_), .B(new_n598_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n595_), .A2(new_n596_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n534_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT72), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n602_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n606_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT73), .B(KEYINPUT74), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT36), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n607_), .A2(new_n618_), .A3(new_n612_), .A4(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT76), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n592_), .B(new_n620_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n622_), .B(new_n623_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n627_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n629_), .A2(new_n592_), .A3(new_n620_), .A4(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n591_), .A2(new_n450_), .A3(new_n396_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n633_), .A2(KEYINPUT101), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n629_), .A2(new_n620_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n591_), .A2(new_n396_), .A3(new_n636_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n634_), .A2(new_n633_), .B1(new_n637_), .B2(G1gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n633_), .B2(new_n634_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT102), .ZN(G1324gat));
  INV_X1    g440(.A(new_n348_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n591_), .A2(new_n451_), .A3(new_n642_), .A4(new_n632_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n465_), .A2(new_n590_), .A3(new_n642_), .A4(new_n636_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G8gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n646_), .B2(KEYINPUT39), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT103), .B(new_n648_), .C1(new_n645_), .C2(G8gat), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n648_), .A3(G8gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT104), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n643_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT40), .B(new_n643_), .C1(new_n650_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1325gat));
  NAND2_X1  g456(.A1(new_n591_), .A2(new_n636_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G15gat), .B1(new_n658_), .B2(new_n365_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT41), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n591_), .A2(new_n632_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n661_), .A2(G15gat), .A3(new_n365_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n658_), .B2(new_n284_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n284_), .A2(G22gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n661_), .B2(new_n666_), .ZN(G1327gat));
  NOR3_X1   g466(.A1(new_n551_), .A2(new_n589_), .A3(new_n463_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n401_), .A2(new_n402_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n411_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n395_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n671_), .A2(new_n419_), .A3(new_n418_), .A4(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n407_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n283_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n365_), .B1(new_n670_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n397_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n628_), .A2(new_n631_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n669_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT43), .B(new_n632_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n668_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n423_), .B2(new_n632_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n678_), .A2(new_n669_), .A3(new_n679_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(KEYINPUT44), .A3(new_n668_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n684_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n398_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n678_), .A2(new_n668_), .A3(new_n629_), .A4(new_n620_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n396_), .A2(new_n554_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT105), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n692_), .B2(new_n694_), .ZN(G1328gat));
  AOI21_X1  g494(.A(new_n558_), .B1(new_n689_), .B2(new_n642_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n692_), .A2(G36gat), .A3(new_n348_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT45), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n696_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  INV_X1    g501(.A(new_n365_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n684_), .A2(G43gat), .A3(new_n703_), .A4(new_n688_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT107), .B(G43gat), .Z(new_n706_));
  OAI21_X1  g505(.A(new_n706_), .B1(new_n692_), .B2(new_n365_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n705_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n705_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n709_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n704_), .A2(new_n707_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT108), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT47), .B1(new_n714_), .B2(new_n708_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1330gat));
  NAND3_X1  g515(.A1(new_n689_), .A2(G50gat), .A3(new_n283_), .ZN(new_n717_));
  INV_X1    g516(.A(G50gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n692_), .B2(new_n284_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1331gat));
  NOR2_X1   g519(.A1(new_n550_), .A2(new_n588_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n465_), .A2(new_n636_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n465_), .A2(KEYINPUT109), .A3(new_n721_), .A4(new_n636_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(new_n437_), .A3(new_n398_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n465_), .A2(new_n721_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n632_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n396_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1332gat));
  NAND3_X1  g531(.A1(new_n730_), .A2(new_n438_), .A3(new_n642_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G64gat), .B1(new_n726_), .B2(new_n348_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT110), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(G64gat), .C1(new_n726_), .C2(new_n348_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n735_), .A2(KEYINPUT48), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT48), .B1(new_n735_), .B2(new_n737_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n733_), .B1(new_n738_), .B2(new_n739_), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n726_), .B2(new_n365_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT49), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n365_), .A2(G71gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n729_), .B2(new_n743_), .ZN(G1334gat));
  OR3_X1    g543(.A1(new_n729_), .A2(G78gat), .A3(new_n284_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G78gat), .B1(new_n726_), .B2(new_n284_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT111), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(G78gat), .C1(new_n726_), .C2(new_n284_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n747_), .A2(KEYINPUT50), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT50), .B1(new_n747_), .B2(new_n749_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n745_), .B1(new_n750_), .B2(new_n751_), .ZN(G1335gat));
  NAND2_X1  g551(.A1(new_n721_), .A2(new_n464_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n423_), .A2(new_n753_), .A3(new_n636_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n396_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n396_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n757_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g557(.A(G92gat), .B1(new_n754_), .B2(new_n642_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n348_), .A2(new_n329_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n756_), .B2(new_n760_), .ZN(G1337gat));
  AOI21_X1  g560(.A(new_n467_), .B1(new_n756_), .B2(new_n703_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n365_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n754_), .B2(new_n763_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n468_), .B1(new_n756_), .B2(new_n283_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770_));
  INV_X1    g569(.A(new_n753_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n283_), .B(new_n771_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G106gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n773_), .B2(KEYINPUT52), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n767_), .A2(KEYINPUT112), .A3(new_n768_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n769_), .A2(new_n774_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n754_), .A2(new_n468_), .A3(new_n283_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(new_n781_), .A3(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n579_), .A2(G229gat), .A3(G233gat), .ZN(new_n785_));
  INV_X1    g584(.A(new_n583_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n569_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n552_), .B1(new_n787_), .B2(new_n572_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT115), .B(new_n789_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n549_), .A2(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n513_), .A2(new_n517_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n497_), .A2(new_n515_), .A3(new_n514_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT68), .B1(new_n534_), .B2(new_n535_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n796_), .A2(new_n797_), .A3(new_n509_), .A4(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT114), .B1(new_n537_), .B2(new_n510_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n537_), .B2(new_n510_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n537_), .A2(new_n510_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n802_), .B(new_n801_), .C1(new_n807_), .C2(new_n804_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n543_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n806_), .A2(new_n811_), .A3(new_n808_), .A4(new_n543_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n810_), .A2(new_n588_), .A3(new_n547_), .A4(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n795_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n814_), .B2(new_n636_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n810_), .A2(new_n794_), .A3(new_n547_), .A4(new_n812_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n679_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT116), .B1(new_n816_), .B2(new_n817_), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n816_), .A2(KEYINPUT116), .A3(new_n817_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n815_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n814_), .A2(KEYINPUT57), .A3(new_n636_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n631_), .A2(new_n628_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n820_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n816_), .A2(KEYINPUT116), .A3(new_n817_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n826_), .B1(new_n830_), .B2(KEYINPUT117), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n463_), .B1(new_n824_), .B2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n550_), .A2(new_n632_), .A3(new_n589_), .A4(new_n463_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT54), .Z(new_n834_));
  OAI21_X1  g633(.A(new_n784_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n825_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n815_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n830_), .B2(KEYINPUT117), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n464_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n833_), .B(KEYINPUT54), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(KEYINPUT118), .A3(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n349_), .A2(new_n365_), .A3(new_n398_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n835_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n588_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n830_), .A2(KEYINPUT119), .A3(new_n837_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n825_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT119), .B1(new_n830_), .B2(new_n837_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n464_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n847_), .B1(new_n851_), .B2(new_n840_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n843_), .B2(KEYINPUT59), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n853_), .A2(new_n588_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n845_), .B1(new_n854_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g654(.A(new_n360_), .B1(new_n550_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n844_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n360_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n853_), .A2(new_n551_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n360_), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n464_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n862_), .B(new_n852_), .C1(new_n843_), .C2(KEYINPUT59), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n835_), .A2(new_n841_), .A3(new_n463_), .A4(new_n842_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n860_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT120), .B1(new_n863_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n853_), .A2(new_n861_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n869_), .A3(new_n865_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n870_), .ZN(G1342gat));
  NOR2_X1   g670(.A1(new_n843_), .A2(new_n636_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n853_), .A2(new_n679_), .ZN(new_n873_));
  MUX2_X1   g672(.A(new_n872_), .B(new_n873_), .S(G134gat), .Z(G1343gat));
  AND3_X1   g673(.A1(new_n835_), .A2(new_n365_), .A3(new_n841_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n284_), .A2(new_n642_), .A3(new_n398_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n588_), .A3(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT121), .B(G141gat), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n877_), .B(new_n878_), .Z(G1344gat));
  NAND3_X1  g678(.A1(new_n875_), .A2(new_n551_), .A3(new_n876_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n875_), .A2(new_n463_), .A3(new_n876_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  NAND2_X1  g683(.A1(new_n875_), .A2(new_n876_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n679_), .A2(G162gat), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n886_), .B(KEYINPUT122), .Z(new_n887_));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n885_), .A2(new_n636_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n222_), .ZN(G1347gat));
  NAND2_X1  g689(.A1(new_n851_), .A2(new_n840_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n365_), .A2(new_n396_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n642_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n283_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n288_), .B1(new_n896_), .B2(new_n588_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n897_), .A2(KEYINPUT62), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n588_), .A3(new_n305_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(KEYINPUT62), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n898_), .A2(new_n899_), .A3(new_n900_), .ZN(G1348gat));
  AOI21_X1  g700(.A(G176gat), .B1(new_n896_), .B2(new_n551_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n835_), .A2(new_n284_), .A3(new_n841_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n835_), .A2(new_n841_), .A3(KEYINPUT123), .A4(new_n284_), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n289_), .B(new_n550_), .C1(new_n905_), .C2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n893_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n902_), .B1(new_n907_), .B2(new_n908_), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n906_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n910_), .A2(new_n463_), .A3(new_n908_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n296_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n464_), .A2(new_n315_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n911_), .A2(new_n912_), .B1(new_n896_), .B2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n895_), .B2(new_n632_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n896_), .A2(new_n316_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n636_), .ZN(G1351gat));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n284_), .A2(new_n396_), .A3(new_n348_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n835_), .A2(new_n841_), .A3(new_n365_), .A4(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n589_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n918_), .B1(new_n921_), .B2(G197gat), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(G197gat), .ZN(new_n923_));
  INV_X1    g722(.A(G197gat), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n920_), .A2(KEYINPUT124), .A3(new_n924_), .A4(new_n589_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n922_), .A2(new_n923_), .A3(new_n925_), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n920_), .A2(new_n550_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT125), .B(G204gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1353gat));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930_));
  NAND2_X1  g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n463_), .A2(new_n931_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n875_), .A2(new_n930_), .A3(new_n919_), .A4(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  INV_X1    g733(.A(new_n932_), .ZN(new_n935_));
  OAI21_X1  g734(.A(KEYINPUT126), .B1(new_n920_), .B2(new_n935_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n933_), .A2(new_n934_), .A3(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n933_), .B2(new_n936_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1354gat));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n920_), .A2(new_n940_), .A3(new_n632_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n920_), .A2(new_n636_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1355gat));
endmodule


