//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT92), .ZN(new_n211_));
  XOR2_X1   g010(.A(G197gat), .B(G204gat), .Z(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT21), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G204gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(KEYINPUT21), .B(new_n216_), .C1(new_n212_), .C2(KEYINPUT91), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n212_), .A2(KEYINPUT21), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n214_), .A2(new_n217_), .B1(new_n211_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT25), .B(G183gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT86), .B(KEYINPUT23), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(new_n228_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT95), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n232_), .A2(KEYINPUT95), .A3(new_n233_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n227_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G169gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT96), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n222_), .B1(new_n240_), .B2(new_n221_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n228_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n229_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n231_), .B2(new_n242_), .ZN(new_n244_));
  INV_X1    g043(.A(G183gat), .ZN(new_n245_));
  INV_X1    g044(.A(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(KEYINPUT97), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT97), .B1(new_n244_), .B2(new_n247_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n241_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n219_), .A2(new_n238_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT20), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT92), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n210_), .B(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n255_), .B(new_n217_), .C1(KEYINPUT21), .C2(new_n212_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n211_), .A2(new_n218_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n224_), .A2(new_n233_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT25), .B1(new_n260_), .B2(new_n245_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n245_), .A2(KEYINPUT25), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n225_), .B(new_n261_), .C1(new_n262_), .C2(new_n260_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n263_), .A3(new_n244_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n232_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(new_n220_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n264_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n253_), .A2(KEYINPUT102), .B1(new_n258_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT102), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n252_), .A2(new_n270_), .A3(KEYINPUT20), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n209_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n219_), .B1(new_n251_), .B2(new_n238_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT20), .B1(new_n258_), .B2(new_n268_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n208_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n206_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n208_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n208_), .B1(new_n258_), .B2(new_n268_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(new_n252_), .A3(KEYINPUT20), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(new_n206_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT27), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n205_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n282_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n288_), .A2(G228gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(G228gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(G233gat), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT93), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT3), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT2), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(KEYINPUT1), .B2(new_n299_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(KEYINPUT1), .B2(new_n299_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n296_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(new_n294_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n298_), .A2(new_n302_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308_));
  OAI211_X1 g107(.A(KEYINPUT90), .B(new_n293_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n298_), .A2(new_n302_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(new_n306_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(new_n292_), .A3(KEYINPUT29), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n258_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT90), .B1(new_n307_), .B2(new_n308_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n291_), .B1(new_n219_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(KEYINPUT94), .A3(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G78gat), .B(G106gat), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G22gat), .B(G50gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n307_), .A2(new_n323_), .A3(new_n308_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n322_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n326_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n324_), .A3(new_n321_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n318_), .A2(new_n320_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n320_), .B1(new_n318_), .B2(new_n330_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n315_), .A2(new_n317_), .ZN(new_n333_));
  OAI22_X1  g132(.A1(new_n331_), .A2(new_n332_), .B1(KEYINPUT94), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n318_), .A2(new_n330_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n319_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n333_), .A2(KEYINPUT94), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n318_), .A2(new_n320_), .A3(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n287_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342_));
  XOR2_X1   g141(.A(G113gat), .B(G120gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT98), .B1(new_n307_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n312_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n312_), .A2(new_n346_), .A3(KEYINPUT98), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT4), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT99), .B1(new_n347_), .B2(KEYINPUT4), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT99), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n312_), .A2(new_n346_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n351_), .A2(new_n353_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G85gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT0), .B(G57gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n359_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G15gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n268_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G71gat), .B(G99gat), .ZN(new_n375_));
  INV_X1    g174(.A(G43gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n374_), .B(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n380_), .A2(KEYINPUT88), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n344_), .B(KEYINPUT31), .Z(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n380_), .B2(KEYINPUT88), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n382_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n341_), .A2(new_n371_), .A3(new_n386_), .ZN(new_n387_));
  AND4_X1   g186(.A1(new_n371_), .A2(new_n284_), .A3(new_n340_), .A4(new_n286_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT33), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n350_), .A2(KEYINPUT4), .B1(new_n354_), .B2(new_n357_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n360_), .B1(new_n390_), .B2(new_n353_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n391_), .B2(new_n366_), .ZN(new_n392_));
  AND4_X1   g191(.A1(new_n389_), .A2(new_n359_), .A3(new_n366_), .A4(new_n361_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(new_n352_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT100), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n350_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n350_), .A2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n353_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n395_), .B(new_n367_), .C1(new_n397_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n280_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n205_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n285_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT101), .B1(new_n394_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n369_), .A2(KEYINPUT33), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n391_), .A2(new_n389_), .A3(new_n366_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT101), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n281_), .A2(new_n285_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n400_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n401_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n272_), .A2(new_n275_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n370_), .B(new_n413_), .C1(new_n412_), .C2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n405_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n340_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n388_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n387_), .B1(new_n418_), .B2(new_n386_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT103), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G29gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G43gat), .B(G50gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n421_), .B(new_n422_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n424_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT15), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G15gat), .B(G22gat), .ZN(new_n432_));
  INV_X1    g231(.A(G1gat), .ZN(new_n433_));
  INV_X1    g232(.A(G8gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G1gat), .B(G8gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OR3_X1    g238(.A1(new_n431_), .A2(KEYINPUT82), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT82), .B1(new_n431_), .B2(new_n439_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n429_), .A2(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G229gat), .A2(G233gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n429_), .B(new_n439_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n444_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n442_), .A2(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G113gat), .B(G141gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT83), .ZN(new_n451_));
  XOR2_X1   g250(.A(G169gat), .B(G197gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n449_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT84), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n449_), .A2(new_n453_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n449_), .A2(new_n453_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n419_), .A2(new_n420_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n420_), .B1(new_n419_), .B2(new_n460_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  XOR2_X1   g263(.A(G85gat), .B(G92gat), .Z(new_n465_));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(KEYINPUT67), .ZN(new_n469_));
  INV_X1    g268(.A(G99gat), .ZN(new_n470_));
  INV_X1    g269(.A(G106gat), .ZN(new_n471_));
  OAI22_X1  g270(.A1(new_n467_), .A2(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(KEYINPUT67), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n474_));
  AND2_X1   g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n464_), .B(new_n465_), .C1(new_n477_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n479_), .A2(new_n483_), .A3(new_n480_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n475_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n472_), .A2(KEYINPUT68), .A3(new_n476_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n486_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(KEYINPUT70), .A3(new_n465_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT8), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT70), .B1(new_n492_), .B2(new_n465_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n482_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n477_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT66), .B(G85gat), .ZN(new_n498_));
  INV_X1    g297(.A(G92gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(KEYINPUT9), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n465_), .A2(KEYINPUT9), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT65), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n497_), .B(new_n501_), .C1(new_n503_), .C2(G106gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G57gat), .B(G64gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT11), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G71gat), .B(G78gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n508_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n505_), .A2(KEYINPUT11), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n496_), .A2(new_n504_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n496_), .B2(new_n504_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT12), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT64), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n496_), .A2(new_n504_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n513_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT71), .ZN(new_n523_));
  INV_X1    g322(.A(new_n518_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n516_), .A2(new_n521_), .A3(new_n526_), .A4(new_n518_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G120gat), .B(G148gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(G176gat), .B(G204gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n523_), .A2(new_n525_), .A3(new_n527_), .A4(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n534_), .A2(KEYINPUT13), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT13), .B1(new_n534_), .B2(new_n536_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT73), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n438_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(new_n513_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT17), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT79), .ZN(new_n545_));
  NOR2_X1   g344(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n546_));
  AND2_X1   g345(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n544_), .B(new_n545_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G127gat), .B(G155gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT81), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT17), .B1(new_n545_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n543_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n548_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n544_), .A2(new_n554_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n520_), .A2(new_n429_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n431_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n496_), .A2(new_n504_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n568_), .A2(KEYINPUT35), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n562_), .A2(new_n565_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT35), .A3(new_n568_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(KEYINPUT35), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n562_), .A2(new_n572_), .A3(new_n565_), .A4(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT77), .ZN(new_n576_));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT36), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n571_), .A2(new_n581_), .A3(new_n578_), .A4(new_n573_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n579_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT78), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT37), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n583_), .B(new_n587_), .ZN(new_n588_));
  NOR4_X1   g387(.A1(new_n463_), .A2(new_n540_), .A3(new_n561_), .A4(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n433_), .A3(new_n370_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT38), .ZN(new_n591_));
  INV_X1    g390(.A(new_n419_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n580_), .A2(new_n582_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n539_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n454_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(new_n560_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT104), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n371_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n591_), .B1(new_n433_), .B2(new_n602_), .ZN(G1324gat));
  INV_X1    g402(.A(new_n287_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G8gat), .B1(new_n598_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT39), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n589_), .A2(new_n434_), .A3(new_n287_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g408(.A(new_n386_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(G15gat), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n611_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n589_), .A2(new_n616_), .A3(new_n386_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT106), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT106), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n614_), .A2(new_n617_), .A3(new_n621_), .A4(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(G1326gat));
  INV_X1    g422(.A(G22gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n600_), .A2(new_n601_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(new_n340_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT42), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n589_), .A2(new_n624_), .A3(new_n340_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1327gat));
  NOR2_X1   g428(.A1(new_n583_), .A2(new_n560_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n539_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n419_), .A2(new_n460_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT103), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n419_), .A2(new_n420_), .A3(new_n460_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n631_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G29gat), .B1(new_n635_), .B2(new_n370_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n419_), .A2(new_n588_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n560_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n419_), .A2(KEYINPUT43), .A3(new_n588_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n639_), .A2(KEYINPUT44), .A3(new_n597_), .A4(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(new_n597_), .A3(new_n640_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n370_), .A2(G29gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n636_), .B1(new_n647_), .B2(new_n648_), .ZN(G1328gat));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n604_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n641_), .A2(new_n642_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n641_), .A2(new_n642_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n604_), .A2(G36gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT108), .B1(new_n635_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n631_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n658_), .B(new_n656_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n655_), .B1(new_n657_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n635_), .A2(KEYINPUT108), .A3(new_n656_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n660_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(KEYINPUT45), .ZN(new_n665_));
  AOI22_X1  g464(.A1(new_n654_), .A2(G36gat), .B1(new_n662_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n650_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n662_), .A2(new_n665_), .ZN(new_n669_));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n643_), .B2(new_n651_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT109), .B(KEYINPUT46), .C1(new_n669_), .C2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n668_), .A2(new_n672_), .ZN(G1329gat));
  NAND4_X1  g472(.A1(new_n643_), .A2(G43gat), .A3(new_n386_), .A4(new_n646_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n635_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n376_), .B1(new_n675_), .B2(new_n610_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n635_), .B2(new_n340_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n340_), .A2(G50gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n647_), .B2(new_n680_), .ZN(G1331gat));
  XNOR2_X1  g480(.A(new_n593_), .B(new_n587_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n595_), .A2(new_n560_), .A3(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT110), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n592_), .A2(new_n454_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(KEYINPUT110), .B2(new_n683_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G57gat), .B1(new_n687_), .B2(new_n370_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT111), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n455_), .A2(new_n560_), .A3(new_n459_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n592_), .A2(new_n593_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n540_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(G57gat), .A3(new_n370_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n689_), .A2(new_n694_), .ZN(G1332gat));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n687_), .A2(new_n696_), .A3(new_n287_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n693_), .A2(new_n287_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(G64gat), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT48), .B(new_n696_), .C1(new_n693_), .C2(new_n287_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT112), .Z(G1333gat));
  OAI21_X1  g502(.A(G71gat), .B1(new_n692_), .B2(new_n610_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(G71gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n687_), .A2(new_n707_), .A3(new_n386_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1334gat));
  OAI21_X1  g508(.A(G78gat), .B1(new_n692_), .B2(new_n417_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT50), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n417_), .A2(G78gat), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT114), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n687_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1335gat));
  AND3_X1   g514(.A1(new_n540_), .A2(new_n685_), .A3(new_n630_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G85gat), .B1(new_n716_), .B2(new_n370_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n639_), .A2(new_n640_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n539_), .A2(new_n454_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n370_), .A2(new_n498_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT115), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n717_), .B1(new_n721_), .B2(new_n723_), .ZN(G1336gat));
  OAI21_X1  g523(.A(G92gat), .B1(new_n720_), .B2(new_n604_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n716_), .A2(new_n499_), .A3(new_n287_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1337gat));
  AOI21_X1  g526(.A(new_n470_), .B1(new_n721_), .B2(new_n386_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n610_), .A2(new_n503_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n716_), .B2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n718_), .A2(new_n340_), .A3(new_n719_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G106gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT52), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n737_), .A3(G106gat), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n716_), .A2(new_n471_), .A3(new_n340_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1339gat));
  INV_X1    g544(.A(KEYINPUT59), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n341_), .A2(new_n370_), .A3(new_n386_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT123), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n523_), .A2(new_n749_), .A3(new_n527_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n513_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n564_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n496_), .A2(new_n504_), .A3(new_n513_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n519_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT12), .B1(new_n564_), .B2(new_n751_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n524_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n516_), .A2(new_n521_), .A3(KEYINPUT55), .A4(new_n518_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n750_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n533_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT56), .ZN(new_n761_));
  AOI211_X1 g560(.A(new_n761_), .B(new_n535_), .C1(new_n750_), .C2(new_n758_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n454_), .B(new_n536_), .C1(new_n760_), .C2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n534_), .A2(new_n536_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n442_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n453_), .B1(new_n447_), .B2(new_n444_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n449_), .A2(new_n453_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n763_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT57), .B1(new_n769_), .B2(new_n583_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n771_), .B(new_n593_), .C1(new_n763_), .C2(new_n768_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT119), .B1(new_n536_), .B2(new_n767_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n536_), .A2(KEYINPUT119), .A3(new_n767_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n760_), .A2(new_n762_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n682_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n759_), .A2(new_n533_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n761_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n533_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n774_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n536_), .A2(KEYINPUT119), .A3(new_n767_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n780_), .A2(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT121), .B1(new_n784_), .B2(KEYINPUT58), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n776_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n778_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n560_), .B1(new_n773_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n690_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n690_), .A2(new_n791_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n588_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n539_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n794_), .B2(new_n539_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n746_), .B(new_n748_), .C1(new_n790_), .C2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT122), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n789_), .A2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT122), .B(new_n778_), .C1(new_n785_), .C2(new_n788_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n773_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n798_), .B1(new_n803_), .B2(new_n561_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n748_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n460_), .B(new_n799_), .C1(new_n806_), .C2(new_n746_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G113gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n454_), .A2(new_n536_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n768_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n583_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n771_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n769_), .A2(KEYINPUT57), .A3(new_n583_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n800_), .B2(new_n789_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n560_), .B1(new_n816_), .B2(new_n802_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n748_), .B1(new_n817_), .B2(new_n798_), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n818_), .A2(G113gat), .A3(new_n596_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n808_), .A2(new_n819_), .ZN(G1340gat));
  OAI211_X1 g619(.A(new_n540_), .B(new_n799_), .C1(new_n806_), .C2(new_n746_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G120gat), .ZN(new_n822_));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n539_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n806_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(G1341gat));
  OAI211_X1 g625(.A(new_n560_), .B(new_n799_), .C1(new_n806_), .C2(new_n746_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G127gat), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n818_), .A2(G127gat), .A3(new_n561_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1342gat));
  INV_X1    g629(.A(KEYINPUT124), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n804_), .A2(new_n583_), .A3(new_n805_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(G134gat), .ZN(new_n833_));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT124), .B(new_n834_), .C1(new_n818_), .C2(new_n583_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n799_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n818_), .B2(KEYINPUT59), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n682_), .A2(new_n834_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n833_), .A2(new_n835_), .B1(new_n837_), .B2(new_n838_), .ZN(G1343gat));
  NOR2_X1   g638(.A1(new_n386_), .A2(new_n417_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n370_), .A3(new_n604_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(KEYINPUT125), .Z(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n803_), .A2(new_n561_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n796_), .A2(new_n797_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n454_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n540_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT126), .B(G148gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1345gat));
  NAND2_X1  g650(.A1(new_n846_), .A2(new_n560_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1346gat));
  INV_X1    g653(.A(KEYINPUT127), .ZN(new_n855_));
  INV_X1    g654(.A(G162gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n846_), .B2(new_n588_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n804_), .A2(G162gat), .A3(new_n583_), .A4(new_n843_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n583_), .A2(G162gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n846_), .A2(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n804_), .A2(new_n682_), .A3(new_n843_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n861_), .B(KEYINPUT127), .C1(new_n862_), .C2(new_n856_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n859_), .A2(new_n863_), .ZN(G1347gat));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n610_), .A2(new_n604_), .A3(new_n370_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n417_), .B(new_n866_), .C1(new_n790_), .C2(new_n798_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n865_), .B(G169gat), .C1(new_n867_), .C2(new_n596_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n773_), .A2(new_n789_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n561_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n340_), .B1(new_n871_), .B2(new_n845_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n454_), .A3(new_n866_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n865_), .B1(new_n873_), .B2(G169gat), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n872_), .A2(new_n240_), .A3(new_n454_), .A4(new_n866_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n869_), .B1(new_n874_), .B2(new_n875_), .ZN(G1348gat));
  NAND3_X1  g675(.A1(new_n872_), .A2(new_n595_), .A3(new_n866_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n804_), .A2(new_n340_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n540_), .A2(G176gat), .A3(new_n866_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n877_), .A2(new_n221_), .B1(new_n878_), .B2(new_n879_), .ZN(G1349gat));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n560_), .A3(new_n866_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n866_), .A2(new_n560_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n226_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n881_), .A2(new_n245_), .B1(new_n872_), .B2(new_n883_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n867_), .B2(new_n682_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n593_), .A2(new_n225_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n867_), .B2(new_n886_), .ZN(G1351gat));
  NAND3_X1  g686(.A1(new_n840_), .A2(new_n371_), .A3(new_n287_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n804_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n454_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n540_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  NAND2_X1  g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  AND4_X1   g694(.A1(new_n560_), .A2(new_n889_), .A3(new_n894_), .A4(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n889_), .B2(new_n560_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1354gat));
  INV_X1    g697(.A(new_n889_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G218gat), .B1(new_n899_), .B2(new_n682_), .ZN(new_n900_));
  INV_X1    g699(.A(G218gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n889_), .A2(new_n901_), .A3(new_n593_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1355gat));
endmodule


