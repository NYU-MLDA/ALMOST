//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n965_, new_n966_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n975_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT81), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G43gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT79), .B(G176gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(KEYINPUT22), .B(G169gat), .Z(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(KEYINPUT78), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT22), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(G169gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(KEYINPUT80), .A3(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT79), .B(G176gat), .Z(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n215_), .B(new_n213_), .C1(new_n211_), .C2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT23), .ZN(new_n221_));
  OR2_X1    g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n221_), .A2(new_n222_), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(new_n219_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n227_), .A2(KEYINPUT24), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n221_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(KEYINPUT24), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT77), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n229_), .B(new_n231_), .C1(new_n235_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n224_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n207_), .B1(new_n241_), .B2(KEYINPUT82), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n244_), .A3(new_n207_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G127gat), .ZN(new_n249_));
  INV_X1    g048(.A(G134gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G127gat), .A2(G134gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G113gat), .ZN(new_n254_));
  INV_X1    g053(.A(G113gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n255_), .A3(new_n252_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n254_), .A2(G120gat), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(G120gat), .B1(new_n254_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT31), .Z(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT83), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n248_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n246_), .A2(new_n261_), .A3(new_n247_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT28), .B(G106gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G22gat), .B(G50gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G228gat), .A2(G233gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT84), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n274_), .B(new_n275_), .C1(new_n272_), .C2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n271_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n276_), .A2(new_n272_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n275_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n286_), .A2(KEYINPUT85), .A3(new_n281_), .A4(new_n274_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n272_), .B(KEYINPUT3), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT86), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT2), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(KEYINPUT2), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n288_), .B(new_n293_), .C1(new_n292_), .C2(new_n290_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n278_), .A2(new_n280_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n283_), .A2(new_n287_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT89), .B(KEYINPUT29), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G211gat), .B(G218gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT21), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n301_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n300_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n299_), .A2(new_n301_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n296_), .A2(new_n298_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G197gat), .B(G204gat), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n303_), .A3(new_n300_), .ZN(new_n310_));
  OR3_X1    g109(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n310_), .A2(KEYINPUT87), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT87), .B1(new_n310_), .B2(new_n311_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n270_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n287_), .A2(new_n283_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n294_), .A2(new_n295_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT29), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT87), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n306_), .B2(new_n302_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n310_), .A2(KEYINPUT87), .A3(new_n311_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n269_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT88), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  AOI221_X4 g126(.A(new_n268_), .B1(new_n270_), .B2(new_n307_), .C1(new_n320_), .C2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n320_), .A2(new_n327_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n307_), .A2(new_n270_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n267_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n266_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n315_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n324_), .A2(new_n326_), .A3(KEYINPUT88), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n330_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n268_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n329_), .A2(new_n330_), .A3(new_n267_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n266_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n296_), .A2(new_n325_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT90), .B(G78gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n332_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n332_), .B2(new_n339_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT91), .Z(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT19), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n350_));
  NAND2_X1  g149(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n350_), .A2(new_n227_), .A3(new_n230_), .A4(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n221_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n351_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n353_), .A2(KEYINPUT93), .A3(new_n234_), .A4(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n355_), .A2(new_n234_), .A3(new_n221_), .A4(new_n352_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n215_), .A2(new_n216_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n356_), .A2(new_n359_), .B1(new_n223_), .B2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n306_), .A2(new_n302_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT20), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n312_), .A2(new_n313_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(new_n239_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n349_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT18), .B(G64gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G92gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n239_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n361_), .A2(new_n362_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(KEYINPUT20), .A4(new_n348_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n366_), .A2(new_n370_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n366_), .B2(new_n373_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n259_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n318_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n296_), .A2(new_n259_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(KEYINPUT4), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n296_), .A2(new_n259_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n318_), .A2(new_n377_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT94), .B1(new_n387_), .B2(new_n381_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT94), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n378_), .A2(new_n379_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n385_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n386_), .A2(new_n392_), .A3(KEYINPUT33), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G85gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(G1gat), .B(G29gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n384_), .A2(new_n391_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n391_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(KEYINPUT33), .A3(new_n397_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n385_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n405_), .A2(KEYINPUT33), .A3(new_n401_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n376_), .A2(new_n399_), .A3(new_n404_), .A4(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n405_), .A2(new_n401_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT96), .B1(new_n408_), .B2(new_n398_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT96), .ZN(new_n410_));
  NOR4_X1   g209(.A1(new_n405_), .A2(new_n410_), .A3(new_n401_), .A4(new_n397_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n398_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n348_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n223_), .A2(new_n360_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n362_), .A2(new_n416_), .A3(new_n357_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n371_), .A2(KEYINPUT20), .A3(new_n349_), .A4(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n366_), .A2(new_n373_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n414_), .B(KEYINPUT95), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n414_), .A2(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n407_), .B1(new_n413_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n345_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n370_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n366_), .A2(new_n370_), .A3(new_n373_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT27), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n415_), .A2(new_n425_), .A3(new_n418_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n427_), .A2(new_n429_), .A3(KEYINPUT27), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n413_), .B(new_n431_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n265_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n332_), .A2(new_n339_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n342_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n332_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n265_), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n428_), .A2(new_n430_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n410_), .B1(new_n403_), .B2(new_n397_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n411_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n441_), .B(new_n442_), .C1(new_n408_), .C2(new_n398_), .ZN(new_n443_));
  NOR4_X1   g242(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .A4(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n433_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G50gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G29gat), .B(G36gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G43gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n447_), .A2(G43gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n446_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G29gat), .B(G36gat), .Z(new_n452_));
  INV_X1    g251(.A(G43gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(G50gat), .A3(new_n448_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT10), .B(G99gat), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n460_), .B(new_n461_), .C1(new_n462_), .C2(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT64), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(G85gat), .B2(G92gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(G85gat), .B2(G92gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT66), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G85gat), .ZN(new_n470_));
  INV_X1    g269(.A(G92gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT65), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT9), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(KEYINPUT64), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n469_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n469_), .B2(new_n478_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n464_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n482_));
  INV_X1    g281(.A(G99gat), .ZN(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n460_), .A3(new_n461_), .A4(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n474_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n470_), .A2(new_n471_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT67), .B1(new_n491_), .B2(new_n473_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n487_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT8), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n487_), .B(new_n495_), .C1(new_n490_), .C2(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n457_), .A2(new_n481_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G232gat), .A2(G233gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT70), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT34), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n494_), .A2(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n481_), .A2(KEYINPUT69), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n468_), .B2(new_n473_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT66), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n476_), .B1(new_n472_), .B2(new_n477_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n469_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n463_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n504_), .B1(new_n505_), .B2(new_n514_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n449_), .A2(new_n446_), .A3(new_n450_), .ZN(new_n516_));
  AOI21_X1  g315(.A(G50gat), .B1(new_n454_), .B2(new_n448_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT15), .B1(new_n451_), .B2(new_n455_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n498_), .B(new_n503_), .C1(new_n515_), .C2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n501_), .A2(new_n502_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G190gat), .B(G218gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(new_n250_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G162gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n512_), .A2(new_n513_), .ZN(new_n530_));
  AOI211_X1 g329(.A(KEYINPUT69), .B(new_n463_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n497_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n456_), .A2(new_n518_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n451_), .A2(KEYINPUT15), .A3(new_n455_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n523_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n503_), .A4(new_n498_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n524_), .A2(new_n529_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT71), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n524_), .A2(new_n538_), .A3(new_n541_), .A4(new_n529_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n527_), .B(new_n528_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n524_), .B2(new_n538_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT72), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n545_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT72), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(KEYINPUT37), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n554_));
  AOI211_X1 g353(.A(KEYINPUT72), .B(new_n545_), .C1(new_n540_), .C2(new_n542_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n445_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(G57gat), .ZN(new_n559_));
  INV_X1    g358(.A(G64gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G57gat), .A2(G64gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n564_));
  XOR2_X1   g363(.A(G71gat), .B(G78gat), .Z(new_n565_));
  OR2_X1    g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT11), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n567_), .A3(new_n562_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n481_), .A2(new_n570_), .A3(new_n497_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n481_), .B2(new_n497_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(new_n572_), .B2(KEYINPUT12), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n532_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n570_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n504_), .B2(new_n512_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT68), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n571_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n575_), .ZN(new_n584_));
  OAI211_X1 g383(.A(KEYINPUT68), .B(new_n580_), .C1(new_n504_), .C2(new_n512_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n579_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588_));
  INV_X1    g387(.A(G204gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT5), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n226_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT13), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n579_), .A2(new_n586_), .A3(new_n592_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT13), .B1(new_n593_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(G1gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT73), .B(G8gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT14), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G15gat), .B(G22gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n602_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT14), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n607_), .A3(new_n602_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G8gat), .B1(new_n606_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n606_), .A2(new_n609_), .A3(G8gat), .ZN(new_n612_));
  OAI22_X1  g411(.A1(new_n519_), .A2(new_n520_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n606_), .A2(G8gat), .A3(new_n609_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n457_), .A2(new_n615_), .A3(new_n610_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT75), .ZN(new_n618_));
  INV_X1    g417(.A(new_n614_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n457_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n611_), .A2(new_n456_), .A3(new_n612_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT75), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n613_), .A2(new_n623_), .A3(new_n614_), .A4(new_n616_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n618_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G169gat), .B(G197gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT76), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(G113gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(G141gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(new_n630_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n618_), .A2(new_n622_), .A3(new_n624_), .A4(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT74), .B1(new_n615_), .B2(new_n610_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n615_), .A2(KEYINPUT74), .A3(new_n610_), .ZN(new_n637_));
  INV_X1    g436(.A(G231gat), .ZN(new_n638_));
  INV_X1    g437(.A(G233gat), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n636_), .B(new_n637_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n639_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT74), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n611_), .A2(new_n612_), .A3(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n643_), .B2(new_n635_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n570_), .B1(new_n640_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n570_), .A3(new_n644_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT16), .B(G183gat), .ZN(new_n648_));
  INV_X1    g447(.A(G211gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n646_), .A2(new_n647_), .B1(KEYINPUT17), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n647_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n652_), .B(KEYINPUT17), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n655_), .A2(new_n645_), .A3(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n601_), .A2(new_n634_), .A3(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n558_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n602_), .A3(new_n443_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT38), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n445_), .A2(new_n549_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n659_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n413_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1324gat));
  OAI21_X1  g465(.A(G8gat), .B1(new_n664_), .B2(new_n431_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT39), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n660_), .A2(new_n603_), .A3(new_n440_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n664_), .B2(new_n439_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT41), .Z(new_n673_));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n660_), .A2(new_n674_), .A3(new_n265_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1326gat));
  OR2_X1    g475(.A1(new_n345_), .A2(KEYINPUT97), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n345_), .A2(KEYINPUT97), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G22gat), .B1(new_n664_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT42), .ZN(new_n682_));
  INV_X1    g481(.A(G22gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n660_), .A2(new_n683_), .A3(new_n679_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1327gat));
  NOR2_X1   g484(.A1(new_n601_), .A2(new_n634_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n557_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n445_), .A2(new_n687_), .A3(KEYINPUT43), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n438_), .A2(new_n440_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n439_), .A2(new_n443_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n443_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n693_), .A2(new_n431_), .B1(new_n345_), .B2(new_n423_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n694_), .B2(new_n265_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n689_), .B1(new_n695_), .B2(new_n557_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n686_), .B(new_n658_), .C1(new_n688_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n445_), .B2(new_n687_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n695_), .A2(new_n689_), .A3(new_n557_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n702_), .A2(KEYINPUT44), .A3(new_n686_), .A4(new_n658_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n699_), .A2(new_n443_), .A3(new_n703_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(KEYINPUT98), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(KEYINPUT98), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(G29gat), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n658_), .A2(new_n549_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT99), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n686_), .B(new_n710_), .C1(new_n433_), .C2(new_n444_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT100), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n695_), .A2(new_n713_), .A3(new_n686_), .A4(new_n710_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(G29gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n443_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n707_), .A2(new_n717_), .ZN(G1328gat));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n699_), .A2(new_n440_), .A3(new_n703_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n725_));
  INV_X1    g524(.A(G36gat), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n712_), .A2(new_n714_), .A3(new_n726_), .A4(new_n440_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(KEYINPUT101), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(KEYINPUT101), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT101), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n715_), .A2(new_n731_), .A3(new_n726_), .A4(new_n440_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n727_), .A2(KEYINPUT101), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(KEYINPUT45), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n721_), .B(new_n722_), .C1(new_n724_), .C2(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n728_), .A2(new_n729_), .A3(new_n725_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n732_), .B2(new_n733_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n723_), .A2(G36gat), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n739_), .A2(new_n719_), .A3(new_n720_), .A4(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n736_), .A2(new_n741_), .ZN(G1329gat));
  NAND3_X1  g541(.A1(new_n712_), .A2(new_n714_), .A3(new_n265_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n453_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(new_n453_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n439_), .A2(new_n453_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n699_), .A2(new_n703_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT103), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n699_), .A2(new_n751_), .A3(new_n703_), .A4(new_n748_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n747_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n754_), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n756_), .B(new_n747_), .C1(new_n750_), .C2(new_n752_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1330gat));
  NAND3_X1  g557(.A1(new_n715_), .A2(new_n446_), .A3(new_n679_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n699_), .A2(new_n438_), .A3(new_n703_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G50gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1331gat));
  OAI21_X1  g563(.A(new_n634_), .B1(new_n657_), .B2(new_n654_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n600_), .A2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n558_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G57gat), .B1(new_n767_), .B2(new_n443_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n663_), .A2(new_n766_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n769_), .A2(new_n559_), .A3(new_n413_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1332gat));
  OAI21_X1  g570(.A(G64gat), .B1(new_n769_), .B2(new_n431_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT48), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n767_), .A2(new_n560_), .A3(new_n440_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n769_), .B2(new_n439_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT49), .ZN(new_n777_));
  INV_X1    g576(.A(G71gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n767_), .A2(new_n778_), .A3(new_n265_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT107), .Z(G1334gat));
  OAI21_X1  g580(.A(G78gat), .B1(new_n769_), .B2(new_n680_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT50), .ZN(new_n783_));
  INV_X1    g582(.A(G78gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n767_), .A2(new_n784_), .A3(new_n679_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n600_), .A2(new_n633_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n702_), .A2(new_n658_), .A3(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(G85gat), .A3(new_n443_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n695_), .A2(new_n710_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n787_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n470_), .B1(new_n791_), .B2(new_n413_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n789_), .A2(new_n792_), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n788_), .A2(G92gat), .A3(new_n440_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n471_), .B1(new_n791_), .B2(new_n431_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1337gat));
  OR3_X1    g595(.A1(new_n791_), .A2(new_n462_), .A3(new_n439_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n702_), .A2(new_n658_), .A3(new_n265_), .A4(new_n787_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G99gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G99gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g602(.A1(new_n702_), .A2(new_n658_), .A3(new_n438_), .A4(new_n787_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(G106gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n804_), .B2(G106gat), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n438_), .A2(new_n484_), .ZN(new_n808_));
  OAI22_X1  g607(.A1(new_n806_), .A2(new_n807_), .B1(new_n791_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g609(.A(new_n765_), .B1(new_n599_), .B2(new_n597_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n552_), .A2(new_n556_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT109), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n552_), .A2(new_n556_), .A3(new_n811_), .A4(new_n814_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n813_), .A2(KEYINPUT54), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT54), .B1(new_n813_), .B2(new_n815_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n633_), .A2(new_n596_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n820_));
  INV_X1    g619(.A(new_n577_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n505_), .A2(new_n514_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n497_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n823_), .A2(new_n573_), .A3(new_n584_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n824_), .B2(KEYINPUT55), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n579_), .A2(KEYINPUT110), .A3(new_n826_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n823_), .A2(new_n573_), .B1(KEYINPUT111), .B2(new_n575_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n575_), .A2(KEYINPUT111), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n574_), .A2(new_n578_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n575_), .A2(new_n826_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n825_), .A2(new_n827_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n592_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n833_), .A2(KEYINPUT56), .A3(new_n834_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n819_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n533_), .A2(new_n534_), .B1(new_n615_), .B2(new_n610_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n621_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n613_), .A2(KEYINPUT112), .A3(new_n616_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n619_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n614_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n630_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n632_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT57), .B(new_n547_), .C1(new_n839_), .C2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n819_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n833_), .A2(KEYINPUT56), .A3(new_n834_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n834_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n848_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(KEYINPUT115), .A3(KEYINPUT57), .A4(new_n547_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT114), .B1(new_n847_), .B2(new_n598_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n846_), .A2(new_n596_), .A3(new_n860_), .A4(new_n632_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n837_), .A2(new_n838_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(KEYINPUT58), .A3(new_n862_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT37), .B1(new_n548_), .B2(new_n551_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n554_), .A2(new_n555_), .A3(new_n553_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n865_), .B(new_n867_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n851_), .A2(new_n858_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n549_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT113), .B1(new_n872_), .B2(KEYINPUT57), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n848_), .B1(new_n866_), .B2(new_n852_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n874_), .B(new_n875_), .C1(new_n876_), .C2(new_n549_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n658_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n818_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n690_), .A2(new_n443_), .A3(new_n265_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT116), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n884_), .B(new_n881_), .C1(new_n818_), .C2(new_n879_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n255_), .B(new_n633_), .C1(new_n883_), .C2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n881_), .A2(KEYINPUT59), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n875_), .B1(new_n876_), .B2(new_n549_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n851_), .A2(new_n889_), .A3(new_n870_), .A4(new_n858_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n890_), .A2(new_n658_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n813_), .A2(new_n815_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n813_), .A2(KEYINPUT54), .A3(new_n815_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n888_), .B1(new_n891_), .B2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n881_), .B1(new_n818_), .B2(new_n879_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n897_), .B(new_n633_), .C1(new_n898_), .C2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G113gat), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n886_), .A2(new_n887_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n887_), .B1(new_n886_), .B2(new_n901_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1340gat));
  OR2_X1    g703(.A1(new_n883_), .A2(new_n885_), .ZN(new_n905_));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n600_), .B2(KEYINPUT60), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT118), .B1(new_n906_), .B2(KEYINPUT60), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n905_), .B(new_n909_), .C1(new_n910_), .C2(new_n907_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n898_), .A2(new_n899_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n897_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G120gat), .B1(new_n913_), .B2(new_n600_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n914_), .ZN(G1341gat));
  NOR3_X1   g714(.A1(new_n913_), .A2(new_n249_), .A3(new_n658_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n658_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G127gat), .B1(new_n905_), .B2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1342gat));
  NAND2_X1  g718(.A1(new_n905_), .A2(new_n549_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n913_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT119), .B(G134gat), .Z(new_n922_));
  NOR2_X1   g721(.A1(new_n687_), .A2(new_n922_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n920_), .A2(new_n250_), .B1(new_n921_), .B2(new_n923_), .ZN(G1343gat));
  NOR3_X1   g723(.A1(new_n345_), .A2(new_n440_), .A3(new_n265_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n880_), .A2(new_n443_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n880_), .A2(KEYINPUT120), .A3(new_n443_), .A4(new_n925_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n634_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT121), .B(G141gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1344gat));
  AOI21_X1  g731(.A(new_n600_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n933_));
  INV_X1    g732(.A(G148gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1345gat));
  AOI21_X1  g734(.A(new_n658_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n936_));
  XOR2_X1   g735(.A(KEYINPUT61), .B(G155gat), .Z(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT122), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n936_), .B(new_n938_), .ZN(G1346gat));
  NAND2_X1  g738(.A1(new_n928_), .A2(new_n929_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G162gat), .B1(new_n940_), .B2(new_n549_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n687_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(G162gat), .B2(new_n942_), .ZN(G1347gat));
  NAND2_X1  g742(.A1(new_n691_), .A2(new_n440_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n679_), .A2(new_n944_), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n633_), .B(new_n945_), .C1(new_n891_), .C2(new_n896_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n946_), .A2(new_n947_), .A3(G169gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(KEYINPUT123), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n947_), .B1(new_n946_), .B2(G169gat), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n945_), .B1(new_n891_), .B2(new_n896_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n633_), .A2(new_n216_), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n952_), .B(KEYINPUT124), .Z(new_n953_));
  OAI22_X1  g752(.A1(new_n949_), .A2(new_n950_), .B1(new_n951_), .B2(new_n953_), .ZN(G1348gat));
  INV_X1    g753(.A(new_n951_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n208_), .B1(new_n955_), .B2(new_n601_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n944_), .A2(new_n600_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n438_), .B1(new_n818_), .B2(new_n879_), .ZN(new_n958_));
  AND2_X1   g757(.A1(new_n958_), .A2(G176gat), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n956_), .B1(new_n957_), .B2(new_n959_), .ZN(G1349gat));
  NOR3_X1   g759(.A1(new_n951_), .A2(new_n658_), .A3(new_n232_), .ZN(new_n961_));
  INV_X1    g760(.A(G183gat), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n958_), .A2(new_n917_), .A3(new_n440_), .A4(new_n691_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n961_), .B1(new_n962_), .B2(new_n963_), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n951_), .B2(new_n687_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n549_), .A2(new_n233_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n951_), .B2(new_n966_), .ZN(G1351gat));
  NAND2_X1  g766(.A1(new_n693_), .A2(new_n439_), .ZN(new_n968_));
  OR2_X1    g767(.A1(new_n968_), .A2(KEYINPUT125), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n431_), .B1(new_n968_), .B2(KEYINPUT125), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n880_), .A2(new_n969_), .A3(new_n970_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(new_n633_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g773(.A1(new_n971_), .A2(new_n600_), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n975_), .B(new_n589_), .ZN(G1353gat));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977_));
  INV_X1    g776(.A(KEYINPUT63), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n978_), .A2(new_n649_), .ZN(new_n979_));
  INV_X1    g778(.A(new_n979_), .ZN(new_n980_));
  NAND4_X1  g779(.A1(new_n972_), .A2(new_n977_), .A3(new_n917_), .A4(new_n980_), .ZN(new_n981_));
  NAND4_X1  g780(.A1(new_n880_), .A2(new_n917_), .A3(new_n969_), .A4(new_n970_), .ZN(new_n982_));
  OAI21_X1  g781(.A(KEYINPUT126), .B1(new_n982_), .B2(new_n979_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n981_), .A2(new_n983_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n978_), .A2(new_n649_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  NAND4_X1  g785(.A1(new_n981_), .A2(new_n978_), .A3(new_n983_), .A4(new_n649_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n986_), .A2(new_n987_), .ZN(G1354gat));
  AOI21_X1  g787(.A(G218gat), .B1(new_n972_), .B2(new_n549_), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n971_), .A2(new_n687_), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n989_), .B1(G218gat), .B2(new_n990_), .ZN(G1355gat));
endmodule


