//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n958_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n204_), .B1(G155gat), .B2(G162gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(G155gat), .A3(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT89), .ZN(new_n207_));
  AOI22_X1  g006(.A1(new_n203_), .A2(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n204_), .A2(KEYINPUT89), .A3(G155gat), .A4(G162gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n202_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(new_n203_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  INV_X1    g013(.A(G141gat), .ZN(new_n215_));
  INV_X1    g014(.A(G148gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n213_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT90), .B1(new_n210_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n203_), .B1(new_n211_), .B2(KEYINPUT1), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n207_), .B1(new_n203_), .B2(KEYINPUT1), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n209_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n202_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n217_), .A2(new_n233_), .A3(new_n220_), .A4(new_n218_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(new_n203_), .A3(new_n212_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G127gat), .B(G134gat), .Z(new_n238_));
  XOR2_X1   g037(.A(G113gat), .B(G120gat), .Z(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  NAND3_X1  g039(.A1(new_n225_), .A2(new_n237_), .A3(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n210_), .A2(new_n224_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n238_), .B(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G1gat), .B(G29gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G85gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT0), .B(G57gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  AND3_X1   g049(.A1(new_n241_), .A2(KEYINPUT4), .A3(new_n244_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n225_), .A2(new_n252_), .A3(new_n237_), .A4(new_n240_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n246_), .B(new_n250_), .C1(new_n251_), .C2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n253_), .A2(new_n254_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n241_), .A2(KEYINPUT4), .A3(new_n244_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n243_), .A2(new_n230_), .A3(new_n235_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n230_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n236_), .B1(new_n230_), .B2(new_n235_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n259_), .B1(new_n262_), .B2(new_n240_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n257_), .A2(new_n258_), .B1(new_n263_), .B2(new_n245_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n256_), .B(KEYINPUT101), .C1(new_n264_), .C2(new_n250_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n246_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n250_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT101), .B1(new_n269_), .B2(new_n256_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(G15gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT30), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT22), .B(G169gat), .ZN(new_n279_));
  INV_X1    g078(.A(G176gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT85), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(KEYINPUT85), .A3(new_n280_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n278_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT86), .B1(new_n286_), .B2(KEYINPUT23), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT86), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(G183gat), .A4(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(KEYINPUT84), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n294_), .A3(KEYINPUT23), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT87), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n300_));
  AOI211_X1 g099(.A(new_n300_), .B(new_n297_), .C1(new_n291_), .C2(new_n295_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n285_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(new_n294_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n289_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n286_), .A2(KEYINPUT23), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G169gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(new_n280_), .A3(KEYINPUT83), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT83), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(G169gat), .B2(G176gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT24), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n308_), .A2(new_n310_), .A3(KEYINPUT24), .A4(new_n277_), .ZN(new_n314_));
  INV_X1    g113(.A(G183gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT25), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G183gat), .ZN(new_n318_));
  INV_X1    g117(.A(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT26), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT26), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G190gat), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n316_), .A2(new_n318_), .A3(new_n320_), .A4(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n306_), .A2(new_n313_), .A3(new_n314_), .A4(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G71gat), .B(G99gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G43gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n302_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n302_), .B2(new_n324_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n276_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT31), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n302_), .A2(new_n324_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n275_), .A3(new_n327_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n330_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n331_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n243_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n335_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n275_), .B1(new_n334_), .B2(new_n327_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT31), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n240_), .B1(new_n342_), .B2(new_n336_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n271_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G228gat), .A2(G233gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT92), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT21), .ZN(new_n348_));
  INV_X1    g147(.A(G218gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G211gat), .ZN(new_n350_));
  INV_X1    g149(.A(G211gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G218gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n350_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G197gat), .B(G204gat), .Z(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n348_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G197gat), .B(G204gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT95), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(KEYINPUT95), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n356_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  OAI221_X1 g163(.A(KEYINPUT21), .B1(new_n357_), .B2(new_n358_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n225_), .A2(KEYINPUT29), .A3(new_n237_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n347_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n242_), .A2(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n371_), .A2(new_n366_), .A3(new_n346_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n262_), .B2(KEYINPUT29), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376_));
  INV_X1    g175(.A(new_n374_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n376_), .B(new_n377_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  OAI211_X1 g182(.A(new_n378_), .B(new_n375_), .C1(new_n369_), .C2(new_n372_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n380_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(G8gat), .B(G36gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT19), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n312_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n314_), .A2(new_n323_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT23), .B1(new_n292_), .B2(new_n294_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n305_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n298_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n400_), .A2(new_n296_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n396_), .B1(new_n366_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT100), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n406_), .A2(new_n407_), .B1(new_n332_), .B2(new_n367_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n366_), .A2(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT20), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT100), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n395_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n302_), .A2(new_n366_), .A3(new_n324_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n281_), .A2(new_n277_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n306_), .B2(new_n298_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n296_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT97), .B1(new_n416_), .B2(new_n399_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n323_), .A2(new_n398_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT97), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n296_), .A4(new_n314_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n415_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n413_), .B(KEYINPUT20), .C1(new_n366_), .C2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n422_), .A2(new_n394_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n392_), .B1(new_n412_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n332_), .A2(new_n367_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n395_), .A2(KEYINPUT20), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n421_), .B2(new_n366_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n422_), .A2(new_n394_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n391_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(KEYINPUT27), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT27), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT20), .B1(new_n421_), .B2(new_n366_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n302_), .A2(new_n366_), .A3(new_n324_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n394_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n425_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n434_), .A2(new_n391_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n391_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n387_), .A2(new_n430_), .A3(new_n438_), .ZN(new_n439_));
  OR3_X1    g238(.A1(new_n344_), .A2(new_n439_), .A3(KEYINPUT103), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT103), .B1(new_n344_), .B2(new_n439_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n243_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n342_), .A2(new_n240_), .A3(new_n336_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(KEYINPUT88), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n380_), .A2(new_n384_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n383_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n380_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n436_), .A2(new_n437_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n258_), .A2(new_n254_), .A3(new_n253_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(KEYINPUT33), .A3(new_n246_), .A4(new_n250_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n258_), .A2(new_n245_), .A3(new_n253_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n263_), .A2(new_n254_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n268_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT98), .B1(new_n256_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n256_), .A2(KEYINPUT98), .A3(new_n462_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n454_), .A2(new_n461_), .A3(new_n464_), .A4(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n391_), .A2(KEYINPUT32), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT99), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n269_), .A2(new_n256_), .B1(new_n428_), .B2(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT32), .B(new_n391_), .C1(new_n412_), .C2(new_n423_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n453_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n430_), .A2(new_n438_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT101), .ZN(new_n474_));
  INV_X1    g273(.A(new_n256_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n250_), .B1(new_n455_), .B2(new_n246_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n477_), .B(new_n265_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(KEYINPUT102), .B(new_n448_), .C1(new_n472_), .C2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n271_), .A2(new_n453_), .A3(new_n438_), .A4(new_n430_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n460_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n256_), .A2(KEYINPUT98), .A3(new_n462_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(new_n463_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n483_), .A2(new_n485_), .B1(new_n470_), .B2(new_n469_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n482_), .B1(new_n486_), .B2(new_n453_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT102), .B1(new_n487_), .B2(new_n448_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n442_), .B1(new_n481_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490_));
  INV_X1    g289(.A(G1gat), .ZN(new_n491_));
  INV_X1    g290(.A(G8gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT14), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G1gat), .B(G8gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G29gat), .B(G36gat), .Z(new_n499_));
  XOR2_X1   g298(.A(G43gat), .B(G50gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT80), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n498_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT81), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n496_), .B(new_n497_), .Z(new_n508_));
  INV_X1    g307(.A(new_n502_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n501_), .B(KEYINPUT15), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n498_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n512_), .A3(new_n505_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G169gat), .B(G197gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT82), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n514_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n507_), .A2(new_n519_), .A3(new_n513_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n489_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525_));
  XOR2_X1   g324(.A(G85gat), .B(G92gat), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n529_), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT10), .B(G99gat), .Z(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT6), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n530_), .A2(new_n531_), .A3(new_n534_), .A4(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT8), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n535_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT66), .ZN(new_n541_));
  INV_X1    g340(.A(new_n535_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n539_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT66), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT7), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n541_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n538_), .B1(new_n548_), .B2(new_n526_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n536_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n550_), .A2(new_n538_), .A3(new_n526_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n537_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n553_));
  XOR2_X1   g352(.A(G71gat), .B(G78gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(KEYINPUT11), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT67), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT67), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n554_), .B(new_n558_), .C1(KEYINPUT11), .C2(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n553_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(KEYINPUT68), .A3(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n552_), .A2(KEYINPUT12), .A3(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n563_), .A2(new_n564_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n551_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n547_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n527_), .B1(new_n573_), .B2(new_n541_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n571_), .B1(new_n574_), .B2(new_n538_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n570_), .B1(new_n575_), .B2(new_n537_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n569_), .B1(KEYINPUT12), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n570_), .A3(new_n537_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n525_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n579_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n578_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(new_n576_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n580_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n570_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n552_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT12), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n585_), .A2(new_n589_), .A3(KEYINPUT69), .A4(new_n569_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n581_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G120gat), .B(G148gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n596_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n597_), .A2(new_n598_), .B1(KEYINPUT71), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G134gat), .B(G162gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT76), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n575_), .A2(new_n501_), .A3(new_n537_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n615_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT75), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n618_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n552_), .A2(KEYINPUT74), .A3(new_n511_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT74), .B1(new_n552_), .B2(new_n511_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n619_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n617_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n552_), .A2(new_n511_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n628_), .A2(new_n617_), .A3(new_n619_), .A4(new_n621_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n609_), .B(new_n611_), .C1(new_n627_), .C2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n623_), .A2(new_n624_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n622_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n626_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n616_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n635_), .A2(new_n608_), .A3(new_n607_), .A4(new_n629_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT37), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n508_), .B(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n568_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(new_n567_), .A3(new_n565_), .ZN(new_n644_));
  XOR2_X1   g443(.A(G127gat), .B(G155gat), .Z(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT16), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G183gat), .B(G211gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT17), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n643_), .A2(new_n644_), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT79), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n641_), .B(new_n586_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n648_), .A2(new_n649_), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n653_), .A2(new_n650_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n631_), .A2(KEYINPUT37), .A3(new_n636_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n639_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n604_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n524_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n271_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n491_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT104), .Z(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n664_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT105), .Z(new_n668_));
  AND2_X1   g467(.A1(new_n489_), .A2(new_n637_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n523_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n604_), .A2(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(new_n657_), .A3(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n662_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n666_), .B(new_n668_), .C1(new_n491_), .C2(new_n673_), .ZN(G1324gat));
  AOI21_X1  g473(.A(new_n492_), .B1(new_n672_), .B2(new_n473_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT39), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n661_), .A2(new_n492_), .A3(new_n473_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1325gat));
  INV_X1    g480(.A(new_n448_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n661_), .A2(new_n273_), .A3(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT106), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n273_), .B1(new_n672_), .B2(new_n682_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n687_), .A3(new_n688_), .ZN(G1326gat));
  INV_X1    g488(.A(G22gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n672_), .B2(new_n453_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT42), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n661_), .A2(new_n690_), .A3(new_n453_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1327gat));
  INV_X1    g493(.A(new_n637_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n656_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n604_), .A2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n524_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n662_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n639_), .A2(new_n658_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n489_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n489_), .A2(KEYINPUT107), .A3(new_n701_), .A4(new_n700_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n489_), .A2(new_n701_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT43), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n705_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n671_), .A2(new_n656_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT44), .B1(new_n708_), .B2(new_n710_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n662_), .A2(G29gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n699_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  NAND2_X1  g514(.A1(new_n708_), .A2(new_n710_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n710_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n473_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G36gat), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(G36gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n524_), .A2(new_n697_), .A3(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT45), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(KEYINPUT46), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n722_), .A2(KEYINPUT109), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT109), .B1(new_n722_), .B2(new_n726_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n722_), .A2(new_n725_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n730_));
  OAI22_X1  g529(.A1(new_n727_), .A2(new_n728_), .B1(new_n729_), .B2(new_n730_), .ZN(G1329gat));
  AOI21_X1  g530(.A(G43gat), .B1(new_n698_), .B2(new_n682_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT111), .Z(new_n733_));
  NOR2_X1   g532(.A1(new_n339_), .A2(new_n343_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G43gat), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT110), .B1(new_n713_), .B2(new_n737_), .ZN(new_n738_));
  AND4_X1   g537(.A1(KEYINPUT110), .A2(new_n718_), .A3(new_n719_), .A4(new_n737_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n733_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT47), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n733_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1330gat));
  OAI21_X1  g543(.A(G50gat), .B1(new_n720_), .B2(new_n387_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n387_), .A2(G50gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT112), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n698_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1331gat));
  INV_X1    g548(.A(new_n604_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(new_n659_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n489_), .A2(new_n670_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT113), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(KEYINPUT113), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n662_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  AND4_X1   g557(.A1(new_n670_), .A2(new_n669_), .A3(new_n657_), .A4(new_n604_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n271_), .A2(new_n758_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n757_), .A2(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(G1332gat));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n473_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G64gat), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT48), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n721_), .A2(G64gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n753_), .B2(new_n765_), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n759_), .B2(new_n682_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT49), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n754_), .A2(new_n767_), .A3(new_n682_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT114), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n769_), .A2(new_n773_), .A3(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1334gat));
  INV_X1    g574(.A(G78gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n759_), .B2(new_n453_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT50), .Z(new_n778_));
  NOR2_X1   g577(.A1(new_n387_), .A2(G78gat), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT115), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n753_), .B2(new_n780_), .ZN(G1335gat));
  NOR3_X1   g580(.A1(new_n750_), .A2(new_n523_), .A3(new_n657_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n708_), .A2(new_n782_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT116), .Z(new_n784_));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n271_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n752_), .A2(new_n656_), .A3(new_n695_), .A4(new_n604_), .ZN(new_n786_));
  OR3_X1    g585(.A1(new_n786_), .A2(G85gat), .A3(new_n271_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1336gat));
  OAI21_X1  g587(.A(G92gat), .B1(new_n784_), .B2(new_n721_), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n786_), .A2(G92gat), .A3(new_n721_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1337gat));
  INV_X1    g590(.A(new_n786_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n792_), .A2(new_n735_), .A3(new_n532_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n783_), .A2(new_n682_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G99gat), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n533_), .A3(new_n453_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n783_), .A2(new_n453_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G106gat), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT52), .B(new_n533_), .C1(new_n783_), .C2(new_n453_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT53), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n797_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1339gat));
  AND2_X1   g605(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n807_));
  NOR4_X1   g606(.A1(new_n604_), .A2(new_n659_), .A3(new_n523_), .A4(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n660_), .A2(new_n670_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n808_), .B1(new_n809_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  INV_X1    g613(.A(new_n596_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n581_), .A2(new_n816_), .A3(new_n590_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n552_), .A2(KEYINPUT12), .A3(new_n568_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT12), .B1(new_n552_), .B2(new_n586_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n580_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n569_), .B(new_n578_), .C1(KEYINPUT12), .C2(new_n576_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n820_), .A2(KEYINPUT55), .B1(new_n582_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n815_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n823_), .A2(KEYINPUT56), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n817_), .A2(new_n822_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n815_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT118), .ZN(new_n829_));
  INV_X1    g628(.A(new_n827_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n824_), .A2(new_n829_), .A3(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n523_), .A2(new_n597_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n504_), .A2(new_n505_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n510_), .A2(new_n512_), .A3(new_n506_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n518_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n514_), .A2(new_n517_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n834_), .A2(new_n835_), .B1(new_n599_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n637_), .A2(KEYINPUT57), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n814_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI22_X1  g642(.A1(new_n832_), .A2(new_n831_), .B1(new_n823_), .B2(KEYINPUT56), .ZN(new_n844_));
  INV_X1    g643(.A(new_n833_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n835_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n599_), .A2(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n842_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(KEYINPUT120), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n843_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n824_), .A2(new_n828_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n840_), .A2(new_n597_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(KEYINPUT58), .A3(new_n853_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n701_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n695_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(KEYINPUT57), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT119), .B(new_n862_), .C1(new_n841_), .C2(new_n695_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n851_), .A2(new_n858_), .A3(new_n861_), .A4(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n813_), .B1(new_n864_), .B2(new_n656_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n439_), .A2(new_n734_), .A3(new_n271_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n813_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n862_), .B1(new_n841_), .B2(new_n695_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT120), .B1(new_n848_), .B2(new_n849_), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n814_), .B(new_n842_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n870_), .B(new_n858_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n869_), .B1(new_n874_), .B2(new_n657_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n867_), .A2(KEYINPUT59), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n868_), .A2(new_n877_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT122), .B(G113gat), .Z(new_n879_));
  NOR2_X1   g678(.A1(new_n670_), .A2(new_n879_), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT123), .Z(new_n881_));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n858_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n861_), .A2(new_n863_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n656_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n869_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(KEYINPUT121), .A3(new_n866_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n883_), .A2(new_n888_), .A3(new_n523_), .ZN(new_n889_));
  INV_X1    g688(.A(G113gat), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n878_), .A2(new_n881_), .B1(new_n889_), .B2(new_n890_), .ZN(G1340gat));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n887_), .B2(new_n866_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n813_), .B1(new_n656_), .B2(new_n873_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n876_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n604_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT124), .B1(new_n893_), .B2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n750_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n868_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n897_), .A2(G120gat), .A3(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n750_), .A2(KEYINPUT60), .ZN(new_n902_));
  MUX2_X1   g701(.A(new_n902_), .B(KEYINPUT60), .S(G120gat), .Z(new_n903_));
  NAND3_X1  g702(.A1(new_n883_), .A2(new_n888_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(G1341gat));
  INV_X1    g704(.A(G127gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n657_), .B2(KEYINPUT125), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(KEYINPUT125), .B2(new_n906_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n883_), .A2(new_n888_), .A3(new_n657_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n878_), .A2(new_n908_), .B1(new_n909_), .B2(new_n906_), .ZN(G1342gat));
  NAND3_X1  g709(.A1(new_n868_), .A2(new_n701_), .A3(new_n877_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(G134gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n883_), .A2(new_n888_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n637_), .A2(G134gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1343gat));
  NAND3_X1  g714(.A1(new_n721_), .A2(new_n662_), .A3(new_n453_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n865_), .A2(new_n682_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n523_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n604_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n657_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1346gat));
  INV_X1    g723(.A(G162gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n917_), .A2(new_n925_), .A3(new_n695_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n917_), .A2(new_n701_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n925_), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n875_), .A2(new_n387_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n721_), .A2(new_n662_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n682_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n523_), .A2(new_n279_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT127), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n931_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n875_), .A2(new_n523_), .A3(new_n387_), .A4(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n937_), .A2(G169gat), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n937_), .B2(G169gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n935_), .B1(new_n939_), .B2(new_n940_), .ZN(G1348gat));
  NAND2_X1  g740(.A1(new_n932_), .A2(new_n604_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n865_), .A2(new_n453_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n750_), .A2(new_n280_), .A3(new_n931_), .ZN(new_n944_));
  AOI22_X1  g743(.A1(new_n942_), .A2(new_n280_), .B1(new_n943_), .B2(new_n944_), .ZN(G1349gat));
  NOR2_X1   g744(.A1(new_n931_), .A2(new_n656_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  AOI211_X1 g746(.A(new_n947_), .B(new_n929_), .C1(new_n316_), .C2(new_n318_), .ZN(new_n948_));
  AOI21_X1  g747(.A(G183gat), .B1(new_n943_), .B2(new_n946_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1350gat));
  NAND4_X1  g749(.A1(new_n932_), .A2(new_n320_), .A3(new_n322_), .A4(new_n695_), .ZN(new_n951_));
  AND2_X1   g750(.A1(new_n932_), .A2(new_n701_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(new_n319_), .ZN(G1351gat));
  NAND3_X1  g752(.A1(new_n473_), .A2(new_n271_), .A3(new_n453_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n865_), .A2(new_n682_), .A3(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n523_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g756(.A1(new_n955_), .A2(new_n604_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g758(.A(KEYINPUT63), .B(G211gat), .C1(new_n955_), .C2(new_n657_), .ZN(new_n960_));
  XOR2_X1   g759(.A(KEYINPUT63), .B(G211gat), .Z(new_n961_));
  AND3_X1   g760(.A1(new_n955_), .A2(new_n657_), .A3(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n960_), .A2(new_n962_), .ZN(G1354gat));
  NAND3_X1  g762(.A1(new_n955_), .A2(new_n349_), .A3(new_n695_), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n955_), .A2(new_n701_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n964_), .B1(new_n965_), .B2(new_n349_), .ZN(G1355gat));
endmodule


