//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT73), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT74), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G134gat), .B(G162gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT36), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n206_), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT67), .B(KEYINPUT6), .Z(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n216_), .B(new_n217_), .C1(new_n218_), .C2(KEYINPUT68), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT7), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n218_), .A2(new_n216_), .A3(new_n217_), .A4(KEYINPUT68), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n213_), .A2(new_n215_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n213_), .A2(new_n215_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(G85gat), .ZN(new_n231_));
  INV_X1    g030(.A(G92gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(KEYINPUT9), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n224_), .A2(KEYINPUT9), .A3(new_n225_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT66), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n238_), .A3(new_n235_), .ZN(new_n239_));
  OR2_X1    g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n217_), .A3(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n230_), .A2(new_n237_), .A3(new_n239_), .A4(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n223_), .A2(KEYINPUT8), .A3(new_n226_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n229_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G29gat), .B(G36gat), .Z(new_n246_));
  XOR2_X1   g045(.A(G43gat), .B(G50gat), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT15), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n245_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n252_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n229_), .A2(new_n243_), .A3(new_n256_), .A4(new_n244_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G232gat), .A2(G233gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT34), .Z(new_n259_));
  INV_X1    g058(.A(KEYINPUT35), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(new_n257_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT76), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n255_), .A2(new_n257_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n261_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n260_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n263_), .B1(new_n264_), .B2(new_n269_), .ZN(new_n270_));
  AOI211_X1 g069(.A(KEYINPUT76), .B(new_n268_), .C1(new_n255_), .C2(new_n257_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n210_), .B(new_n262_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT78), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n202_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n262_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n239_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n213_), .A2(new_n215_), .A3(new_n242_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n278_), .A2(new_n237_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n253_), .B1(new_n279_), .B2(new_n244_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n257_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n269_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT76), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n264_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n275_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n208_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT77), .B1(new_n210_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n207_), .A2(new_n209_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT36), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT77), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n272_), .B1(new_n285_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n274_), .A2(new_n294_), .ZN(new_n295_));
  OAI221_X1 g094(.A(new_n272_), .B1(new_n273_), .B2(new_n202_), .C1(new_n285_), .C2(new_n293_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G57gat), .B(G64gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT11), .ZN(new_n299_));
  XOR2_X1   g098(.A(G71gat), .B(G78gat), .Z(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n298_), .A2(KEYINPUT11), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n300_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G231gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G15gat), .A2(G22gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(G15gat), .A2(G22gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT79), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n311_), .A2(new_n310_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n309_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G1gat), .B(G8gat), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n313_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n306_), .B(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G127gat), .B(G155gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT16), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G183gat), .B(G211gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT17), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT81), .Z(new_n330_));
  XOR2_X1   g129(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n331_));
  OR3_X1    g130(.A1(new_n323_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n297_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n334_), .B(KEYINPUT82), .Z(new_n335_));
  XNOR2_X1  g134(.A(G120gat), .B(G148gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT5), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G176gat), .B(G204gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n340_), .A2(KEYINPUT71), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n229_), .A2(new_n243_), .A3(new_n304_), .A4(new_n244_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G230gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT64), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT70), .ZN(new_n347_));
  INV_X1    g146(.A(new_n304_), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n349_));
  NAND3_X1  g148(.A1(new_n245_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n304_), .B1(new_n279_), .B2(new_n244_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT12), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(KEYINPUT69), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n350_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n347_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n345_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n343_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n351_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n342_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n356_), .A2(new_n359_), .A3(new_n342_), .ZN(new_n362_));
  AND2_X1   g161(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n361_), .B(new_n362_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n362_), .ZN(new_n366_));
  OAI22_X1  g165(.A1(new_n366_), .A2(new_n360_), .B1(KEYINPUT72), .B2(KEYINPUT13), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n335_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT18), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  AND2_X1   g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G197gat), .ZN(new_n381_));
  INV_X1    g180(.A(G204gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G197gat), .A2(G204gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(KEYINPUT21), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G211gat), .B(G218gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G218gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G211gat), .ZN(new_n389_));
  INV_X1    g188(.A(G211gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G218gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n392_), .A2(KEYINPUT21), .A3(new_n383_), .A4(new_n384_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n387_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G169gat), .ZN(new_n396_));
  AND3_X1   g195(.A1(KEYINPUT90), .A2(G183gat), .A3(G190gat), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT90), .B1(G183gat), .B2(G190gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT23), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(KEYINPUT87), .A2(G183gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(KEYINPUT87), .A2(G183gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n405_), .A2(G190gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n396_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT23), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT23), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n405_), .B2(KEYINPUT25), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G190gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n417_), .A2(new_n415_), .A3(G190gat), .ZN(new_n418_));
  INV_X1    g217(.A(G190gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT88), .B1(new_n419_), .B2(KEYINPUT26), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n412_), .B1(new_n414_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n423_));
  INV_X1    g222(.A(G169gat), .ZN(new_n424_));
  INV_X1    g223(.A(G176gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT89), .B1(G169gat), .B2(G176gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n426_), .A2(KEYINPUT24), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n426_), .A2(new_n427_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(KEYINPUT24), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n394_), .B(new_n407_), .C1(new_n422_), .C2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT20), .ZN(new_n433_));
  INV_X1    g232(.A(new_n394_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT101), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n412_), .B2(new_n437_), .ZN(new_n438_));
  AOI211_X1 g237(.A(KEYINPUT101), .B(new_n436_), .C1(new_n409_), .C2(new_n411_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n396_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n410_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(KEYINPUT90), .A2(G183gat), .A3(G190gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n400_), .B1(new_n444_), .B2(KEYINPUT23), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(new_n426_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n426_), .A2(new_n427_), .ZN(new_n448_));
  AND2_X1   g247(.A1(KEYINPUT99), .A2(KEYINPUT24), .ZN(new_n449_));
  NOR2_X1   g248(.A1(KEYINPUT99), .A2(KEYINPUT24), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT25), .B(G183gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT26), .B(G190gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n445_), .A2(new_n447_), .A3(new_n452_), .A4(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT100), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n448_), .A2(new_n451_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT100), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n447_), .A4(new_n445_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n440_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n433_), .B1(new_n434_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT19), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT98), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT102), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n457_), .A2(new_n460_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n396_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n411_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n444_), .B2(new_n408_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT101), .B1(new_n471_), .B2(new_n436_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n412_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n434_), .B1(new_n468_), .B2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n432_), .A2(KEYINPUT20), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT102), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n465_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n467_), .A2(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n440_), .A2(new_n394_), .A3(new_n457_), .A4(new_n460_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n407_), .B1(new_n422_), .B2(new_n431_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n434_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n484_), .A3(new_n464_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n376_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  AOI211_X1 g286(.A(new_n375_), .B(new_n487_), .C1(new_n467_), .C2(new_n479_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n371_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n477_), .B2(new_n465_), .ZN(new_n490_));
  AOI211_X1 g289(.A(KEYINPUT102), .B(new_n466_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n376_), .B(new_n485_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n440_), .A2(new_n394_), .A3(new_n456_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n484_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n464_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(new_n477_), .B2(new_n465_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n371_), .B1(new_n497_), .B2(new_n375_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n492_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT104), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT104), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n492_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n489_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G155gat), .A2(G162gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G155gat), .A2(G162gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(G141gat), .A2(G148gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT3), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT3), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(KEYINPUT91), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n509_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G141gat), .A2(G148gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT2), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT2), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n514_), .A2(KEYINPUT92), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(G141gat), .A2(G148gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n512_), .A2(KEYINPUT91), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n510_), .A2(KEYINPUT3), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT92), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT93), .B1(new_n509_), .B2(new_n512_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n525_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n522_), .A2(new_n523_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n508_), .B1(new_n518_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n519_), .A2(new_n515_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n506_), .B1(KEYINPUT1), .B2(new_n504_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n504_), .A2(KEYINPUT1), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT29), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n434_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(G228gat), .A3(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n528_), .B2(new_n532_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT91), .B(KEYINPUT3), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT92), .B1(new_n539_), .B2(new_n519_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n516_), .A2(new_n517_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n523_), .B(new_n509_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n524_), .A2(new_n526_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n507_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n532_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(KEYINPUT94), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n538_), .A2(KEYINPUT29), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n394_), .B1(G228gat), .B2(G233gat), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n548_), .A2(KEYINPUT97), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT97), .B1(new_n548_), .B2(new_n549_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n536_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G78gat), .B(G106gat), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT94), .B1(new_n545_), .B2(new_n546_), .ZN(new_n555_));
  AOI211_X1 g354(.A(new_n537_), .B(new_n532_), .C1(new_n544_), .C2(new_n507_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n534_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT96), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G22gat), .B(G50gat), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n559_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n534_), .B(new_n563_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n560_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n553_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n568_), .B(new_n536_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n554_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n554_), .B2(new_n569_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G71gat), .B(G99gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G43gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n483_), .B(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G127gat), .B(G134gat), .Z(new_n576_));
  XOR2_X1   g375(.A(G113gat), .B(G120gat), .Z(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n575_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G227gat), .A2(G233gat), .ZN(new_n580_));
  INV_X1    g379(.A(G15gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT30), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT31), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n579_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n538_), .A2(new_n547_), .A3(new_n578_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n578_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n533_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(KEYINPUT4), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G225gat), .A2(G233gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT4), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n538_), .A2(new_n593_), .A3(new_n547_), .A4(new_n578_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G1gat), .B(G29gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(G85gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT0), .B(G57gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n587_), .A2(KEYINPUT4), .A3(new_n589_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n594_), .A2(new_n592_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n596_), .B(new_n601_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n586_), .A2(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n503_), .A2(new_n572_), .A3(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n595_), .A2(KEYINPUT33), .A3(new_n596_), .A4(new_n601_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n590_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n587_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n602_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n614_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n606_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n606_), .B2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n376_), .A2(KEYINPUT32), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n603_), .A2(new_n606_), .B1(new_n622_), .B2(new_n497_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n480_), .A2(new_n621_), .A3(new_n485_), .ZN(new_n624_));
  AOI22_X1  g423(.A1(new_n615_), .A2(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n548_), .A2(new_n549_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n548_), .A2(KEYINPUT97), .A3(new_n549_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n568_), .B1(new_n630_), .B2(new_n536_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n569_), .ZN(new_n632_));
  OAI22_X1  g431(.A1(new_n631_), .A2(new_n632_), .B1(new_n566_), .B2(new_n565_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n554_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n607_), .A3(new_n634_), .ZN(new_n635_));
  OAI22_X1  g434(.A1(new_n625_), .A2(new_n572_), .B1(new_n635_), .B2(new_n503_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n609_), .B1(new_n636_), .B2(new_n585_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT86), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G169gat), .B(G197gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n639_), .B(new_n640_), .Z(new_n641_));
  NAND2_X1  g440(.A1(new_n256_), .A2(KEYINPUT83), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT83), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n252_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n321_), .A3(new_n320_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n322_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT84), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT84), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n652_), .B(new_n649_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n253_), .A2(new_n322_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT85), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n646_), .A2(new_n649_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n641_), .B1(new_n654_), .B2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n659_), .B(new_n641_), .C1(new_n651_), .C2(new_n653_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n638_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n641_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(KEYINPUT86), .A3(new_n661_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n637_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n370_), .A2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT105), .Z(new_n672_));
  INV_X1    g471(.A(new_n607_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n307_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT38), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n294_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n637_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n369_), .A2(new_n669_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n333_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n680_), .B2(new_n607_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n674_), .A2(new_n675_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n676_), .A2(new_n681_), .A3(new_n682_), .ZN(G1324gat));
  NAND3_X1  g482(.A1(new_n672_), .A2(new_n308_), .A3(new_n503_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n503_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G8gat), .B1(new_n680_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT39), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n688_), .B(new_n690_), .ZN(G1325gat));
  NAND3_X1  g490(.A1(new_n672_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n693_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G15gat), .B1(new_n680_), .B2(new_n585_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT41), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n694_), .A2(new_n695_), .A3(new_n697_), .ZN(G1326gat));
  INV_X1    g497(.A(new_n572_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(G22gat), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT108), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n672_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G22gat), .B1(new_n680_), .B2(new_n699_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT42), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1327gat));
  NAND2_X1  g504(.A1(new_n330_), .A2(new_n332_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n677_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n670_), .A2(new_n368_), .A3(new_n708_), .ZN(new_n709_));
  OR3_X1    g508(.A1(new_n709_), .A2(G29gat), .A3(new_n607_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n295_), .A2(KEYINPUT109), .A3(new_n296_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(KEYINPUT43), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(new_n637_), .B2(new_n297_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n486_), .A2(new_n488_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n614_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n619_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n606_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .A4(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n623_), .A2(new_n624_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n572_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n503_), .A2(new_n635_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n585_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n609_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n297_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n712_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n713_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n679_), .A2(new_n706_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n728_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n732_), .B(new_n729_), .C1(new_n713_), .C2(new_n727_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n673_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n735_), .A2(KEYINPUT110), .A3(G29gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT110), .B1(new_n735_), .B2(G29gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n710_), .B1(new_n736_), .B2(new_n737_), .ZN(G1328gat));
  AOI21_X1  g537(.A(new_n726_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n297_), .B(new_n712_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n730_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n732_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n728_), .A2(KEYINPUT44), .A3(new_n730_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n503_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT111), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n742_), .A2(new_n746_), .A3(new_n503_), .A4(new_n743_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(G36gat), .A3(new_n747_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n709_), .A2(G36gat), .A3(new_n685_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n748_), .A2(new_n751_), .B1(KEYINPUT112), .B2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n746_), .B1(new_n734_), .B2(new_n503_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n747_), .A2(G36gat), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT112), .B(new_n751_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT113), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(G1329gat));
  NOR3_X1   g558(.A1(new_n709_), .A2(G43gat), .A3(new_n585_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n734_), .A2(new_n586_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(G43gat), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g562(.A1(new_n731_), .A2(new_n733_), .A3(new_n699_), .ZN(new_n764_));
  INV_X1    g563(.A(G50gat), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n572_), .A2(new_n765_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT114), .Z(new_n767_));
  OAI22_X1  g566(.A1(new_n764_), .A2(new_n765_), .B1(new_n709_), .B2(new_n767_), .ZN(G1331gat));
  NOR2_X1   g567(.A1(KEYINPUT116), .A2(G57gat), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n668_), .A2(new_n706_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n678_), .A2(new_n369_), .A3(new_n770_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n607_), .A2(KEYINPUT116), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n769_), .B(new_n771_), .C1(G57gat), .C2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n335_), .A2(new_n368_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n637_), .A2(new_n668_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n777_), .A2(KEYINPUT115), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(KEYINPUT115), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n673_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(G57gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n773_), .B1(new_n780_), .B2(new_n781_), .ZN(G1332gat));
  OAI21_X1  g581(.A(G64gat), .B1(new_n771_), .B2(new_n685_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT48), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n685_), .A2(G64gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n776_), .B2(new_n785_), .ZN(G1333gat));
  OAI21_X1  g585(.A(G71gat), .B1(new_n771_), .B2(new_n585_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT49), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n585_), .A2(G71gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n776_), .B2(new_n789_), .ZN(G1334gat));
  OAI21_X1  g589(.A(G78gat), .B1(new_n771_), .B2(new_n699_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT50), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n699_), .A2(G78gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n776_), .B2(new_n793_), .ZN(G1335gat));
  NOR2_X1   g593(.A1(new_n368_), .A2(new_n707_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n775_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(G85gat), .B1(new_n797_), .B2(new_n673_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n739_), .A2(new_n740_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n368_), .A2(new_n668_), .A3(new_n333_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n673_), .A2(new_n231_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n798_), .B1(new_n802_), .B2(new_n803_), .ZN(G1336gat));
  NAND3_X1  g603(.A1(new_n797_), .A2(new_n232_), .A3(new_n503_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n799_), .A2(new_n685_), .A3(new_n801_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n232_), .ZN(G1337gat));
  AOI21_X1  g606(.A(new_n216_), .B1(new_n802_), .B2(new_n586_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n586_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n797_), .B2(new_n809_), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT51), .Z(G1338gat));
  NOR3_X1   g610(.A1(new_n796_), .A2(G106gat), .A3(new_n699_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n802_), .A2(new_n572_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G106gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT52), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n816_), .A3(G106gat), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n819_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n812_), .B(new_n821_), .C1(new_n815_), .C2(new_n817_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1339gat));
  OAI21_X1  g622(.A(new_n357_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n346_), .A2(KEYINPUT70), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT70), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n831_), .B2(new_n354_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n347_), .A2(KEYINPUT55), .A3(new_n355_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT120), .B(new_n357_), .C1(new_n354_), .C2(new_n358_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n826_), .A2(new_n832_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n339_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT56), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n838_), .A3(new_n339_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n356_), .A2(new_n359_), .A3(new_n340_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n837_), .A2(new_n668_), .A3(new_n839_), .A4(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n641_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n843_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n657_), .A2(new_n646_), .A3(new_n650_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n847_), .A2(new_n661_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n366_), .B2(new_n360_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n841_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n294_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(KEYINPUT57), .A3(new_n294_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n837_), .A2(new_n848_), .A3(new_n839_), .A4(new_n840_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n725_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n840_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n836_), .B2(KEYINPUT56), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n861_), .A2(KEYINPUT58), .A3(new_n848_), .A4(new_n839_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n861_), .A2(new_n839_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(KEYINPUT122), .A3(KEYINPUT58), .A4(new_n848_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n859_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n706_), .B1(new_n855_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n869_));
  OR2_X1    g668(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n770_), .A2(new_n368_), .A3(KEYINPUT118), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n297_), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT118), .B1(new_n770_), .B2(new_n368_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n869_), .B(new_n870_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n873_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n869_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n875_), .A2(new_n297_), .A3(new_n876_), .A4(new_n871_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n868_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n607_), .A2(new_n585_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n880_), .A2(new_n699_), .A3(new_n685_), .A4(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(G113gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n884_), .A3(new_n668_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(KEYINPUT59), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n669_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n889_), .B2(new_n884_), .ZN(G1340gat));
  INV_X1    g689(.A(G120gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n368_), .B2(KEYINPUT60), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n883_), .B(new_n892_), .C1(KEYINPUT60), .C2(new_n891_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n368_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n891_), .ZN(G1341gat));
  INV_X1    g694(.A(G127gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n883_), .A2(new_n896_), .A3(new_n333_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n706_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n896_), .ZN(G1342gat));
  INV_X1    g698(.A(G134gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n882_), .B2(new_n294_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n902_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n886_), .A2(new_n888_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n297_), .A2(new_n900_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n903_), .A2(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1343gat));
  NAND4_X1  g706(.A1(new_n685_), .A2(new_n673_), .A3(new_n572_), .A4(new_n585_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n868_), .B2(new_n879_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n668_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n369_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n333_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT61), .B(G155gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  INV_X1    g715(.A(G162gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n909_), .A2(new_n917_), .A3(new_n677_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n909_), .A2(new_n725_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n920_), .B2(new_n917_), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n572_), .A2(new_n608_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT57), .B1(new_n850_), .B2(new_n294_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n852_), .B(new_n677_), .C1(new_n841_), .C2(new_n849_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n297_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n862_), .A2(new_n863_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n862_), .A2(new_n863_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n333_), .B1(new_n925_), .B2(new_n929_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n503_), .B(new_n922_), .C1(new_n930_), .C2(new_n878_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931_), .B2(new_n669_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT62), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(KEYINPUT124), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n880_), .A2(new_n935_), .A3(new_n503_), .A4(new_n922_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT22), .B(G169gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n937_), .A2(new_n668_), .A3(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n933_), .A2(new_n939_), .ZN(G1348gat));
  NAND3_X1  g739(.A1(new_n937_), .A2(new_n425_), .A3(new_n369_), .ZN(new_n941_));
  OAI21_X1  g740(.A(G176gat), .B1(new_n931_), .B2(new_n368_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1349gat));
  OR2_X1    g742(.A1(new_n706_), .A2(new_n453_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n934_), .B2(new_n936_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n931_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n405_), .B1(new_n946_), .B2(new_n333_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948_));
  OR3_X1    g747(.A1(new_n945_), .A2(new_n947_), .A3(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n945_), .B2(new_n947_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n937_), .A2(new_n454_), .A3(new_n677_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n685_), .B1(new_n868_), .B2(new_n879_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n935_), .B1(new_n953_), .B2(new_n922_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n931_), .A2(KEYINPUT124), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n725_), .B1(new_n954_), .B2(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(KEYINPUT126), .B1(new_n956_), .B2(G190gat), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n297_), .B1(new_n934_), .B2(new_n936_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n958_), .A2(new_n959_), .A3(new_n419_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n952_), .B1(new_n957_), .B2(new_n960_), .ZN(G1351gat));
  NAND4_X1  g760(.A1(new_n953_), .A2(new_n607_), .A3(new_n572_), .A4(new_n585_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(new_n669_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT127), .B(G197gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1352gat));
  NOR2_X1   g764(.A1(new_n962_), .A2(new_n368_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(new_n382_), .ZN(G1353gat));
  NOR2_X1   g766(.A1(new_n962_), .A2(new_n706_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n968_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969_));
  XNOR2_X1  g768(.A(KEYINPUT63), .B(G211gat), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n962_), .A2(new_n706_), .A3(new_n970_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n969_), .A2(new_n971_), .ZN(G1354gat));
  OAI21_X1  g771(.A(G218gat), .B1(new_n962_), .B2(new_n297_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n677_), .A2(new_n388_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n962_), .B2(new_n974_), .ZN(G1355gat));
endmodule


