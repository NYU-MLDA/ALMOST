//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G230gat), .A2(G233gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT64), .Z(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT67), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT7), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n218_), .A2(new_n209_), .A3(new_n210_), .A4(KEYINPUT67), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(KEYINPUT68), .A3(new_n224_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n217_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT69), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n212_), .A4(new_n219_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n221_), .A2(new_n223_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n222_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n223_), .A2(KEYINPUT9), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n217_), .A2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(KEYINPUT10), .B(G99gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT65), .B(G106gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n221_), .A2(KEYINPUT9), .A3(new_n223_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT66), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n238_), .A2(new_n245_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n229_), .A2(new_n236_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G57gat), .B(G64gat), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(KEYINPUT11), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(KEYINPUT11), .ZN(new_n251_));
  XOR2_X1   g050(.A(G71gat), .B(G78gat), .Z(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n251_), .A2(new_n252_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n247_), .A2(new_n248_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n244_), .A2(new_n246_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n227_), .A2(new_n228_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(new_n235_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n255_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT70), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n247_), .A2(new_n255_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n208_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n208_), .B1(new_n247_), .B2(new_n255_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n259_), .A2(new_n266_), .A3(new_n260_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n265_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n206_), .B1(new_n264_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n264_), .A2(new_n269_), .A3(new_n206_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT13), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(KEYINPUT13), .A3(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT71), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G127gat), .B(G155gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT16), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G183gat), .B(G211gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G231gat), .A2(G233gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n260_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G1gat), .B(G8gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT79), .ZN(new_n291_));
  OR2_X1    g090(.A1(G15gat), .A2(G22gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G15gat), .A2(G22gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G1gat), .A2(G8gat), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n292_), .A2(new_n293_), .B1(KEYINPUT14), .B2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n291_), .B(new_n295_), .Z(new_n296_));
  NOR2_X1   g095(.A1(new_n260_), .A2(new_n287_), .ZN(new_n297_));
  OR3_X1    g096(.A1(new_n289_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n289_), .B2(new_n297_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT80), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n286_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT17), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT17), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n300_), .B2(new_n286_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G190gat), .B(G218gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G134gat), .B(G162gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n313_));
  XOR2_X1   g112(.A(G29gat), .B(G36gat), .Z(new_n314_));
  XOR2_X1   g113(.A(G43gat), .B(G50gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n313_), .B1(new_n259_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n229_), .A2(new_n236_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(KEYINPUT72), .A3(new_n316_), .A4(new_n257_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G232gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT34), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT35), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT74), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n323_), .A2(KEYINPUT35), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n316_), .B(KEYINPUT15), .ZN(new_n327_));
  AOI211_X1 g126(.A(new_n325_), .B(new_n326_), .C1(new_n259_), .C2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(KEYINPUT74), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n321_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n321_), .B2(new_n328_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n312_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT75), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n321_), .A2(new_n328_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n329_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n321_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n337_));
  XOR2_X1   g136(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n310_), .B(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n343_), .B(new_n312_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n336_), .A2(KEYINPUT77), .A3(new_n337_), .A4(new_n339_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n333_), .A2(new_n342_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT37), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n332_), .A2(new_n340_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT78), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n332_), .A2(new_n340_), .A3(new_n350_), .A4(new_n347_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n346_), .A2(KEYINPUT37), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n281_), .A2(new_n307_), .A3(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G78gat), .B(G106gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT95), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT92), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G211gat), .B(G218gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G197gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G204gat), .ZN(new_n361_));
  INV_X1    g160(.A(G204gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(G197gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(KEYINPUT21), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n360_), .A3(G204gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT21), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n361_), .A2(new_n363_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(KEYINPUT93), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n358_), .B1(new_n364_), .B2(KEYINPUT21), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n365_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G155gat), .ZN(new_n373_));
  INV_X1    g172(.A(G162gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT89), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(G155gat), .B2(G162gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT1), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT90), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n383_), .A3(KEYINPUT1), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n379_), .B2(KEYINPUT1), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n378_), .B(new_n382_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G141gat), .ZN(new_n388_));
  INV_X1    g187(.A(G148gat), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G141gat), .A2(G148gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT2), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n394_), .A2(new_n396_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n380_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n387_), .A2(new_n392_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n357_), .B(new_n372_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT94), .B(new_n372_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n404_));
  AND2_X1   g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n356_), .A2(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n356_), .A3(new_n405_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n355_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n356_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n404_), .A2(new_n405_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n355_), .B(KEYINPUT96), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n407_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n387_), .A2(new_n392_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n399_), .A2(new_n400_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n402_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT28), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT28), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n401_), .A2(new_n420_), .A3(new_n402_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G22gat), .B(G50gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n409_), .A2(new_n415_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n413_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n419_), .A2(new_n421_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n422_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(KEYINPUT91), .A3(new_n423_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n428_), .A2(new_n415_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT97), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n427_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n428_), .A2(new_n415_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n430_), .A2(new_n434_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n409_), .A2(new_n415_), .A3(new_n426_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT97), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G127gat), .B(G134gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(G113gat), .B(G120gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT86), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(G183gat), .A3(G190gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT23), .ZN(new_n451_));
  INV_X1    g250(.A(G183gat), .ZN(new_n452_));
  INV_X1    g251(.A(G190gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT23), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n446_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT88), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n451_), .A2(new_n459_), .A3(new_n454_), .A4(new_n456_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G169gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(G183gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(G183gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n452_), .A2(KEYINPUT25), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n467_), .B1(new_n470_), .B2(new_n465_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT26), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G190gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n453_), .A2(KEYINPUT26), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(KEYINPUT83), .A3(G190gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n464_), .B1(new_n471_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G169gat), .ZN(new_n480_));
  INV_X1    g279(.A(G176gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT24), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G169gat), .A2(G176gat), .ZN(new_n483_));
  OR3_X1    g282(.A1(new_n482_), .A2(KEYINPUT84), .A3(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT84), .B1(new_n482_), .B2(new_n483_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT23), .B1(new_n447_), .B2(new_n449_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n446_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n446_), .A2(KEYINPUT23), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n491_), .B(new_n494_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n479_), .B(new_n486_), .C1(new_n490_), .C2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n463_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G71gat), .B(G99gat), .ZN(new_n498_));
  INV_X1    g297(.A(G43gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n497_), .A2(new_n500_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n445_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n503_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n443_), .B(new_n444_), .Z(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n501_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(G15gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT30), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT31), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n504_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n437_), .A2(new_n442_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n401_), .A2(new_n506_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n392_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n386_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n384_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n375_), .A2(new_n377_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n399_), .A2(new_n400_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n445_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT102), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n517_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n401_), .A2(new_n506_), .A3(KEYINPUT102), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(KEYINPUT4), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G29gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G85gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT0), .B(G57gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n526_), .A2(new_n527_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n532_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n533_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n531_), .B2(new_n540_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n545_), .B2(new_n538_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n532_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n547_));
  NOR4_X1   g346(.A1(new_n547_), .A2(KEYINPUT33), .A3(new_n537_), .A4(new_n544_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n542_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G226gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n372_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n463_), .A2(new_n496_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT99), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(KEYINPUT20), .ZN(new_n557_));
  INV_X1    g356(.A(new_n462_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n487_), .A2(new_n488_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n559_), .A2(new_n489_), .A3(new_n491_), .A4(new_n494_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n560_), .B2(new_n454_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n483_), .B1(new_n482_), .B2(KEYINPUT100), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(KEYINPUT100), .B2(new_n482_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n470_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n473_), .A2(new_n474_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n464_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AND4_X1   g365(.A1(new_n456_), .A2(new_n563_), .A3(new_n451_), .A4(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n372_), .B1(new_n561_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n557_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n556_), .B1(new_n555_), .B2(KEYINPUT20), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n553_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n561_), .A2(new_n372_), .A3(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n497_), .A2(new_n372_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n572_), .A2(KEYINPUT20), .A3(new_n552_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G8gat), .B(G36gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT18), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G64gat), .B(G92gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n571_), .A2(new_n579_), .A3(new_n574_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT101), .A3(new_n582_), .ZN(new_n583_));
  AOI211_X1 g382(.A(KEYINPUT101), .B(new_n579_), .C1(new_n571_), .C2(new_n574_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n549_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n545_), .A2(new_n538_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT103), .ZN(new_n588_));
  NOR4_X1   g387(.A1(new_n547_), .A2(new_n588_), .A3(new_n537_), .A4(new_n544_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n545_), .A2(new_n538_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n588_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n569_), .A2(new_n553_), .A3(new_n570_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n572_), .A2(KEYINPUT20), .A3(new_n573_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n553_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n593_), .A2(KEYINPUT32), .A3(new_n579_), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n579_), .A2(KEYINPUT32), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n575_), .A2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n590_), .A2(new_n592_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n516_), .B1(new_n586_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n590_), .A2(new_n592_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n436_), .B1(new_n427_), .B2(new_n435_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n440_), .A2(KEYINPUT97), .A3(new_n441_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n515_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n515_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT27), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n583_), .A2(new_n585_), .A3(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n593_), .A2(new_n595_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT27), .B(new_n582_), .C1(new_n610_), .C2(new_n579_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n600_), .B1(new_n607_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n291_), .B(new_n295_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n316_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(new_n316_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n327_), .A2(new_n296_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G113gat), .B(G141gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G169gat), .B(G197gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OR3_X1    g426(.A1(new_n623_), .A2(KEYINPUT81), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT81), .B1(new_n623_), .B2(new_n627_), .ZN(new_n629_));
  AOI22_X1  g428(.A1(new_n628_), .A2(new_n629_), .B1(new_n623_), .B2(new_n627_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n613_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n353_), .A2(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n602_), .A2(G1gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n634_), .A2(KEYINPUT38), .A3(new_n635_), .A4(new_n636_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n612_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n515_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n603_), .A2(new_n604_), .A3(new_n515_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n601_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n591_), .A2(KEYINPUT33), .ZN(new_n646_));
  INV_X1    g445(.A(new_n548_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n646_), .A2(new_n647_), .B1(new_n533_), .B2(new_n541_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n582_), .A2(KEYINPUT101), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n579_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n651_), .B2(new_n584_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n596_), .A2(new_n598_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n601_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n641_), .A2(new_n645_), .B1(new_n655_), .B2(new_n516_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n332_), .A2(new_n340_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT105), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n277_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n631_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n307_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n602_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n639_), .A2(new_n640_), .A3(new_n665_), .ZN(G1324gat));
  INV_X1    g465(.A(G8gat), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n634_), .A2(new_n667_), .A3(new_n612_), .A4(new_n635_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n659_), .A2(new_n662_), .A3(new_n612_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n667_), .B1(new_n670_), .B2(KEYINPUT39), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n672_));
  AOI22_X1  g471(.A1(new_n669_), .A2(new_n671_), .B1(KEYINPUT106), .B2(new_n672_), .ZN(new_n673_));
  AND4_X1   g472(.A1(KEYINPUT106), .A2(new_n669_), .A3(new_n672_), .A4(G8gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n668_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n668_), .B(KEYINPUT40), .C1(new_n673_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  NAND2_X1  g478(.A1(new_n663_), .A2(new_n515_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n680_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(new_n680_), .B2(G15gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n515_), .A2(new_n509_), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n681_), .A2(new_n682_), .B1(new_n633_), .B2(new_n683_), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n437_), .A2(new_n442_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n633_), .A2(G22gat), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n685_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n663_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(G22gat), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G22gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n686_), .B1(new_n690_), .B2(new_n691_), .ZN(G1327gat));
  INV_X1    g491(.A(new_n657_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n307_), .A2(new_n693_), .ZN(new_n694_));
  NOR4_X1   g493(.A1(new_n656_), .A2(new_n630_), .A3(new_n277_), .A4(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n601_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n660_), .A2(new_n631_), .A3(new_n307_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n613_), .A2(new_n699_), .A3(new_n352_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n613_), .B2(new_n352_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT44), .B(new_n698_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT108), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n346_), .A2(KEYINPUT37), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n349_), .A2(new_n351_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n656_), .B2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n613_), .A2(new_n699_), .A3(new_n352_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(KEYINPUT44), .A4(new_n698_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n703_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n698_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n601_), .A2(G29gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n696_), .B1(new_n717_), .B2(new_n718_), .ZN(G1328gat));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  INV_X1    g519(.A(G36gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n641_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n712_), .B2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n695_), .A2(new_n721_), .A3(new_n612_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT45), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n695_), .A2(new_n726_), .A3(new_n721_), .A4(new_n612_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n720_), .B1(new_n723_), .B2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n697_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n612_), .B1(new_n731_), .B2(KEYINPUT44), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n703_), .B2(new_n711_), .ZN(new_n733_));
  OAI211_X1 g532(.A(KEYINPUT46), .B(new_n728_), .C1(new_n733_), .C2(new_n721_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1329gat));
  XNOR2_X1  g534(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n515_), .A2(G43gat), .ZN(new_n738_));
  AOI221_X4 g537(.A(new_n738_), .B1(new_n714_), .B2(new_n713_), .C1(new_n703_), .C2(new_n711_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G43gat), .B1(new_n695_), .B2(new_n515_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n740_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n736_), .C1(new_n716_), .C2(new_n738_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1330gat));
  NOR2_X1   g543(.A1(new_n685_), .A2(G50gat), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT111), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n695_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n685_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n712_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G50gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n712_), .B2(new_n749_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n751_), .B2(new_n752_), .ZN(G1331gat));
  NOR3_X1   g552(.A1(new_n352_), .A2(new_n660_), .A3(new_n307_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n613_), .A3(new_n630_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n755_), .A2(KEYINPUT112), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(KEYINPUT112), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n602_), .A2(G57gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n306_), .A2(new_n630_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n659_), .A2(new_n281_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n601_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G57gat), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n759_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT113), .ZN(G1332gat));
  OR3_X1    g564(.A1(new_n755_), .A2(G64gat), .A3(new_n641_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n612_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G64gat), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1333gat));
  OR3_X1    g570(.A1(new_n755_), .A2(G71gat), .A3(new_n642_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n761_), .A2(new_n515_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G71gat), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  OR3_X1    g576(.A1(new_n755_), .A2(G78gat), .A3(new_n685_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n761_), .A2(new_n687_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G78gat), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT50), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT50), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(G1335gat));
  INV_X1    g582(.A(new_n694_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n281_), .A2(new_n613_), .A3(new_n630_), .A4(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(G85gat), .B1(new_n787_), .B2(new_n601_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n789_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n660_), .A2(new_n631_), .A3(new_n306_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n709_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n601_), .A2(G85gat), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT116), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n790_), .A2(new_n791_), .B1(new_n793_), .B2(new_n795_), .ZN(G1336gat));
  AOI21_X1  g595(.A(G92gat), .B1(new_n787_), .B2(new_n612_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n612_), .A2(G92gat), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT117), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n793_), .B2(new_n799_), .ZN(G1337gat));
  AND2_X1   g599(.A1(new_n515_), .A2(new_n239_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n787_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n709_), .A2(new_n515_), .A3(new_n792_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G99gat), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(KEYINPUT118), .A3(KEYINPUT51), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n787_), .A2(new_n801_), .B1(new_n803_), .B2(G99gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n805_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n809_), .B2(new_n808_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n807_), .B1(new_n810_), .B2(new_n812_), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n787_), .A2(new_n687_), .A3(new_n240_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n709_), .A2(new_n687_), .A3(new_n792_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(G106gat), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n815_), .B2(G106gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT53), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n814_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1339gat));
  NOR2_X1   g622(.A1(new_n267_), .A2(new_n268_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n208_), .B1(new_n824_), .B2(new_n262_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n269_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n265_), .B(KEYINPUT55), .C1(new_n267_), .C2(new_n268_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n205_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT56), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n832_), .A3(new_n205_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n831_), .A2(new_n631_), .A3(new_n272_), .A4(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n614_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n627_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n836_), .A2(KEYINPUT120), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n618_), .A2(new_n614_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n836_), .A2(KEYINPUT120), .B1(new_n621_), .B2(new_n838_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n628_), .A2(new_n629_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n273_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n834_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n657_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n272_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n830_), .B2(KEYINPUT56), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n840_), .A3(new_n833_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(KEYINPUT121), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(KEYINPUT121), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n847_), .A2(new_n851_), .A3(new_n840_), .A4(new_n833_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n352_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n842_), .A2(KEYINPUT57), .A3(new_n657_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n845_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n307_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n760_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n706_), .B2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n760_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n352_), .A2(new_n860_), .A3(KEYINPUT54), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n856_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n612_), .A2(new_n602_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n515_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n864_), .A2(new_n685_), .A3(new_n867_), .A4(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n862_), .B1(new_n855_), .B2(new_n307_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n870_), .A2(new_n687_), .A3(new_n866_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n872_));
  OAI211_X1 g671(.A(new_n869_), .B(new_n631_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G113gat), .ZN(new_n874_));
  INV_X1    g673(.A(G113gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(new_n875_), .A3(new_n631_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1340gat));
  OAI211_X1 g676(.A(new_n869_), .B(new_n281_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G120gat), .ZN(new_n879_));
  INV_X1    g678(.A(G120gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n660_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n871_), .B(new_n881_), .C1(KEYINPUT60), .C2(new_n880_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1341gat));
  OAI211_X1 g682(.A(new_n869_), .B(new_n306_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G127gat), .ZN(new_n885_));
  INV_X1    g684(.A(G127gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n871_), .A2(new_n886_), .A3(new_n306_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1342gat));
  INV_X1    g687(.A(new_n658_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n870_), .A2(new_n687_), .A3(new_n889_), .A4(new_n866_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT123), .B1(new_n890_), .B2(G134gat), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT124), .B(G134gat), .Z(new_n892_));
  NOR2_X1   g691(.A1(new_n706_), .A2(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n869_), .B(new_n893_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n864_), .A2(new_n685_), .A3(new_n658_), .A4(new_n867_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  INV_X1    g695(.A(G134gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n891_), .A2(new_n894_), .A3(new_n898_), .ZN(G1343gat));
  NOR2_X1   g698(.A1(new_n870_), .A2(new_n643_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n631_), .A3(new_n865_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n281_), .A3(new_n865_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g703(.A1(new_n900_), .A2(new_n306_), .A3(new_n865_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT61), .B(G155gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1346gat));
  NOR2_X1   g706(.A1(new_n889_), .A2(G162gat), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n864_), .A2(new_n606_), .A3(new_n865_), .A4(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n865_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n870_), .A2(new_n643_), .A3(new_n706_), .A4(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n374_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT125), .B(new_n909_), .C1(new_n911_), .C2(new_n374_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n870_), .A2(new_n687_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n641_), .A2(new_n601_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n515_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n631_), .A3(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT62), .B(G169gat), .C1(new_n921_), .C2(KEYINPUT22), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n870_), .A2(new_n687_), .A3(new_n630_), .A4(new_n919_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT22), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n480_), .B1(new_n924_), .B2(new_n923_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n922_), .B1(new_n926_), .B2(new_n927_), .ZN(G1348gat));
  NAND2_X1  g727(.A1(new_n917_), .A2(new_n920_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n280_), .B2(new_n279_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n277_), .A2(new_n481_), .ZN(new_n931_));
  OAI22_X1  g730(.A1(new_n930_), .A2(new_n481_), .B1(new_n929_), .B2(new_n931_), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n917_), .A2(new_n306_), .A3(new_n920_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n564_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n452_), .B2(new_n933_), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n929_), .B2(new_n706_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n658_), .A2(new_n565_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n929_), .B2(new_n937_), .ZN(G1351gat));
  INV_X1    g737(.A(new_n918_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n870_), .A2(new_n643_), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n631_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n281_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g743(.A(new_n307_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n900_), .A2(new_n918_), .A3(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n947_), .A2(KEYINPUT126), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n946_), .A2(new_n948_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n947_), .B(KEYINPUT126), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n946_), .B2(new_n950_), .ZN(G1354gat));
  NAND2_X1  g750(.A1(new_n940_), .A2(new_n658_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(KEYINPUT127), .ZN(new_n953_));
  NOR4_X1   g752(.A1(new_n870_), .A2(new_n643_), .A3(new_n889_), .A4(new_n939_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955_));
  AOI21_X1  g754(.A(G218gat), .B1(new_n954_), .B2(new_n955_), .ZN(new_n956_));
  AND2_X1   g755(.A1(new_n352_), .A2(G218gat), .ZN(new_n957_));
  AOI22_X1  g756(.A1(new_n953_), .A2(new_n956_), .B1(new_n940_), .B2(new_n957_), .ZN(G1355gat));
endmodule


