//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n965_, new_n966_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_, new_n986_;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT87), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT1), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n203_), .B(new_n206_), .C1(new_n209_), .C2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n207_), .B(KEYINPUT88), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n204_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n203_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n213_), .B(new_n210_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n220_), .A2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n212_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226_));
  INV_X1    g025(.A(G197gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT93), .B1(new_n227_), .B2(G204gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(KEYINPUT21), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n226_), .A2(KEYINPUT21), .ZN(new_n232_));
  XOR2_X1   g031(.A(G197gat), .B(G204gat), .Z(new_n233_));
  NAND4_X1  g032(.A1(new_n233_), .A2(KEYINPUT21), .A3(new_n226_), .A4(new_n228_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G78gat), .B(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n225_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n220_), .A2(new_n221_), .ZN(new_n240_));
  AND3_X1   g039(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n243_), .A2(KEYINPUT89), .A3(new_n218_), .A4(new_n215_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n240_), .A2(new_n244_), .A3(new_n213_), .A4(new_n210_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n239_), .B1(new_n245_), .B2(new_n212_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n236_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT92), .A2(G228gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(G233gat), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n238_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n238_), .B2(new_n248_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n202_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n238_), .A2(new_n248_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n252_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n238_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT94), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G22gat), .B(G50gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT91), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n245_), .A2(new_n265_), .A3(new_n239_), .A4(new_n212_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n261_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n261_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n267_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n256_), .A2(new_n260_), .A3(new_n270_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n273_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT94), .B1(new_n258_), .B2(new_n259_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G120gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(G127gat), .A2(G134gat), .ZN(new_n280_));
  INV_X1    g079(.A(G113gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G127gat), .A2(G134gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n281_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n279_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n285_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(G120gat), .A3(new_n283_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT86), .B(G176gat), .ZN(new_n290_));
  INV_X1    g089(.A(G169gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT22), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT85), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT22), .B(G169gat), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n290_), .B(new_n293_), .C1(new_n294_), .C2(KEYINPUT85), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT83), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G183gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(G190gat), .B1(new_n302_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n297_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n304_), .A3(KEYINPUT25), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT26), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G190gat), .ZN(new_n310_));
  INV_X1    g109(.A(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT26), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT84), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n311_), .A2(KEYINPUT84), .A3(KEYINPUT26), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n307_), .A2(new_n308_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n298_), .A2(new_n299_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(KEYINPUT24), .A3(new_n297_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n296_), .A2(new_n306_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(KEYINPUT30), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n318_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n308_), .A2(new_n307_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n313_), .A2(new_n314_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n303_), .A2(G183gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n301_), .A2(KEYINPUT83), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n311_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n335_), .A2(new_n318_), .B1(G169gat), .B2(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n295_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n327_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n289_), .B1(new_n326_), .B2(new_n338_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n331_), .A2(new_n328_), .B1(new_n336_), .B2(new_n295_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n327_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n325_), .A2(KEYINPUT30), .ZN(new_n342_));
  INV_X1    g141(.A(new_n289_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G15gat), .B(G43gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT31), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n339_), .A2(new_n344_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n339_), .B2(new_n344_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n349_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n339_), .A2(new_n344_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n346_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n353_), .B1(new_n357_), .B2(new_n348_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n278_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT18), .B(G64gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G92gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(new_n320_), .A3(new_n297_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT26), .B(G190gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n322_), .A2(KEYINPUT95), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n322_), .A2(KEYINPUT95), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n319_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n366_), .A2(new_n369_), .A3(new_n372_), .A4(new_n318_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n290_), .A2(new_n294_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n374_), .B(new_n297_), .C1(new_n300_), .C2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n235_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n332_), .A2(new_n337_), .A3(new_n247_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT19), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n378_), .A2(new_n379_), .A3(KEYINPUT20), .A4(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n325_), .B2(new_n235_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n247_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n381_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n364_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n386_), .B(KEYINPUT20), .C1(new_n340_), .C2(new_n247_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n381_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n364_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n382_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(KEYINPUT96), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT96), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n395_), .B(new_n364_), .C1(new_n383_), .C2(new_n387_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT97), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT97), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n399_), .A3(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n343_), .A2(new_n245_), .A3(new_n212_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n224_), .A2(KEYINPUT98), .A3(new_n289_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n245_), .A2(new_n212_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT4), .B1(new_n408_), .B2(KEYINPUT98), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n403_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n405_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(new_n408_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n402_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n410_), .A2(new_n413_), .A3(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n402_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n412_), .A2(new_n403_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n418_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT101), .ZN(new_n426_));
  AND2_X1   g225(.A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n420_), .B1(new_n421_), .B2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n401_), .A2(new_n422_), .A3(new_n426_), .A4(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n378_), .A2(new_n379_), .A3(KEYINPUT20), .A4(new_n390_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(KEYINPUT102), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n389_), .A2(new_n381_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(KEYINPUT102), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT103), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n410_), .A2(new_n413_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n418_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n420_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n435_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(new_n387_), .B2(new_n383_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n360_), .B1(new_n429_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n434_), .A2(new_n392_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(KEYINPUT27), .A3(new_n388_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT27), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n394_), .A2(new_n448_), .A3(new_n396_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n355_), .A2(new_n358_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n278_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n359_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n453_));
  AOI211_X1 g252(.A(new_n450_), .B(new_n441_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n445_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT80), .ZN(new_n456_));
  AND2_X1   g255(.A1(G57gat), .A2(G64gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G57gat), .A2(G64gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT68), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G57gat), .ZN(new_n460_));
  INV_X1    g259(.A(G64gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT68), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G57gat), .A2(G64gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT11), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n468_));
  XOR2_X1   g267(.A(G71gat), .B(G78gat), .Z(new_n469_));
  AND3_X1   g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n466_), .B1(new_n459_), .B2(new_n465_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n470_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n467_), .A2(new_n469_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT69), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n472_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G231gat), .A2(G233gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n473_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n476_), .A2(new_n477_), .A3(new_n472_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(G231gat), .A3(G233gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G1gat), .A2(G8gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT14), .ZN(new_n488_));
  INV_X1    g287(.A(G15gat), .ZN(new_n489_));
  INV_X1    g288(.A(G22gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(G15gat), .A2(G22gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT79), .ZN(new_n494_));
  XOR2_X1   g293(.A(G1gat), .B(G8gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(KEYINPUT79), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n486_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n481_), .A2(new_n500_), .A3(new_n485_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT16), .B(G183gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(G211gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G127gat), .B(G155gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT17), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n504_), .A2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n508_), .A2(KEYINPUT17), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n502_), .A2(new_n513_), .A3(new_n503_), .A4(new_n510_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n456_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n514_), .A3(new_n456_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G190gat), .B(G218gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G134gat), .B(G162gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT76), .B(G29gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G36gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(G43gat), .B(G50gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(G36gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n526_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n529_), .A2(new_n533_), .A3(KEYINPUT15), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT7), .ZN(new_n542_));
  INV_X1    g341(.A(G99gat), .ZN(new_n543_));
  INV_X1    g342(.A(G106gat), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .A4(KEYINPUT67), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT67), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT7), .ZN(new_n547_));
  OAI22_X1  g346(.A1(new_n546_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n541_), .A2(new_n545_), .A3(new_n547_), .A4(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT8), .ZN(new_n550_));
  AND2_X1   g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(G85gat), .A2(G92gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n550_), .B1(new_n549_), .B2(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT70), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(G92gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT65), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT65), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G92gat), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n561_), .A3(G85gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT66), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n552_), .B1(new_n551_), .B2(KEYINPUT9), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT66), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n567_), .A3(new_n563_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT10), .B(G99gat), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n544_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n541_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n549_), .A2(new_n553_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT8), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n554_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n557_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n554_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n578_), .A2(new_n572_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n538_), .A2(new_n577_), .B1(new_n579_), .B2(new_n534_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT34), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(KEYINPUT35), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n580_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n525_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n523_), .B(new_n524_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n583_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT37), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n518_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n455_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  INV_X1    g402(.A(G204gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT5), .ZN(new_n606_));
  INV_X1    g405(.A(G176gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT73), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n608_), .A2(new_n609_), .A3(KEYINPUT74), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT74), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n606_), .B(G176gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n612_), .B2(KEYINPUT73), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n479_), .A2(new_n579_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n578_), .A2(new_n572_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n484_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT64), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT71), .B1(new_n474_), .B2(new_n478_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n482_), .A2(new_n483_), .A3(new_n509_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n622_), .A2(KEYINPUT12), .A3(new_n577_), .A4(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n620_), .B1(new_n479_), .B2(new_n579_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n617_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n614_), .B1(new_n621_), .B2(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n610_), .A2(new_n613_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n621_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n601_), .B(new_n602_), .C1(new_n629_), .C2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n631_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n614_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n630_), .A2(new_n631_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n599_), .A4(new_n600_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n500_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n534_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n494_), .A2(new_n496_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n495_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n646_), .A2(new_n529_), .A3(new_n533_), .A4(new_n497_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n642_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n641_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G113gat), .B(G141gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(new_n291_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(G197gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n643_), .A2(new_n650_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT82), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n643_), .A2(new_n650_), .A3(KEYINPUT82), .A4(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n643_), .A2(new_n650_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n653_), .B(KEYINPUT81), .Z(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n639_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n598_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n441_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n665_), .A2(G1gat), .A3(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT38), .Z(new_n668_));
  NAND2_X1  g467(.A1(new_n429_), .A2(new_n444_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n360_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n452_), .A2(new_n453_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n450_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n666_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n593_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n518_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n664_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G1gat), .B1(new_n679_), .B2(new_n666_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n668_), .A2(new_n680_), .ZN(G1324gat));
  OAI21_X1  g480(.A(G8gat), .B1(new_n679_), .B2(new_n673_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT39), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n665_), .A2(G8gat), .A3(new_n673_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n683_), .A2(KEYINPUT40), .A3(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n679_), .B2(new_n359_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT104), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT104), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n665_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n489_), .A3(new_n451_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n694_), .A2(new_n696_), .A3(new_n697_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n679_), .B2(new_n278_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  INV_X1    g499(.A(new_n278_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(new_n490_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT105), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(new_n705_), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1327gat));
  AND3_X1   g506(.A1(new_n512_), .A2(new_n514_), .A3(new_n456_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n515_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n709_), .A2(new_n633_), .A3(new_n637_), .A4(new_n662_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n589_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n595_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n445_), .B2(new_n454_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT107), .B1(new_n713_), .B2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT43), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n719_), .B(new_n716_), .C1(new_n445_), .C2(new_n454_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n712_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT108), .B1(new_n723_), .B2(KEYINPUT44), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n722_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n712_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n724_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n723_), .A2(KEYINPUT44), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n731_), .A2(G29gat), .A3(new_n441_), .A4(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G29gat), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n455_), .A2(new_n676_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n710_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n737_), .B2(new_n666_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1328gat));
  AOI21_X1  g540(.A(new_n673_), .B1(new_n723_), .B2(KEYINPUT44), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n731_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G36gat), .ZN(new_n744_));
  NAND2_X1  g543(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n745_));
  OR2_X1    g544(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n737_), .A2(G36gat), .A3(new_n673_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT45), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .A4(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n530_), .B1(new_n731_), .B2(new_n742_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT110), .B(KEYINPUT46), .C1(new_n751_), .C2(new_n748_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1329gat));
  NAND4_X1  g552(.A1(new_n731_), .A2(G43gat), .A3(new_n451_), .A4(new_n732_), .ZN(new_n754_));
  INV_X1    g553(.A(G43gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n737_), .B2(new_n359_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g557(.A(new_n737_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G50gat), .B1(new_n759_), .B2(new_n701_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n278_), .B1(new_n724_), .B2(new_n730_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n732_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1331gat));
  AOI22_X1  g562(.A1(new_n656_), .A2(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n638_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n678_), .A2(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n767_), .A2(new_n460_), .A3(new_n666_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n598_), .A2(new_n766_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G57gat), .B1(new_n770_), .B2(new_n441_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n768_), .A2(new_n771_), .ZN(G1332gat));
  OAI21_X1  g571(.A(G64gat), .B1(new_n767_), .B2(new_n673_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT48), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n461_), .A3(new_n450_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1333gat));
  INV_X1    g575(.A(G71gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n770_), .A2(new_n777_), .A3(new_n451_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n677_), .A2(new_n359_), .A3(new_n765_), .ZN(new_n779_));
  OR3_X1    g578(.A1(new_n779_), .A2(KEYINPUT111), .A3(new_n777_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT111), .B1(new_n779_), .B2(new_n777_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(KEYINPUT49), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT49), .B1(new_n780_), .B2(new_n781_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT112), .B(new_n778_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1334gat));
  NAND3_X1  g587(.A1(new_n678_), .A2(new_n701_), .A3(new_n766_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n789_), .A2(G78gat), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n791_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(KEYINPUT50), .A3(new_n793_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n278_), .A2(G78gat), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT114), .Z(new_n799_));
  OAI211_X1 g598(.A(new_n796_), .B(new_n797_), .C1(new_n769_), .C2(new_n799_), .ZN(G1335gat));
  NAND2_X1  g599(.A1(new_n766_), .A2(new_n709_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n735_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G85gat), .B1(new_n804_), .B2(new_n441_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n801_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(new_n666_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n805_), .B1(new_n808_), .B2(G85gat), .ZN(G1336gat));
  NAND4_X1  g608(.A1(new_n806_), .A2(new_n559_), .A3(new_n561_), .A4(new_n450_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n558_), .B1(new_n803_), .B2(new_n673_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1337gat));
  OAI21_X1  g611(.A(G99gat), .B1(new_n807_), .B2(new_n359_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n451_), .A2(new_n570_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n813_), .B(new_n814_), .C1(new_n803_), .C2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n278_), .B(new_n801_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n819_), .B2(new_n544_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n725_), .A2(new_n701_), .A3(new_n802_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(G106gat), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n803_), .A2(G106gat), .A3(new_n278_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n818_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  AOI211_X1 g626(.A(KEYINPUT116), .B(new_n825_), .C1(new_n820_), .C2(new_n823_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n819_), .A2(KEYINPUT52), .A3(new_n544_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n822_), .B1(new_n821_), .B2(G106gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n826_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT116), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n824_), .A2(new_n818_), .A3(new_n826_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT53), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n830_), .A2(new_n836_), .ZN(G1339gat));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n633_), .A2(new_n637_), .A3(new_n764_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n709_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n597_), .A2(new_n839_), .A3(KEYINPUT54), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n662_), .B1(new_n631_), .B2(new_n612_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n624_), .A2(new_n615_), .A3(new_n627_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n620_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n628_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n624_), .A2(new_n625_), .A3(new_n627_), .A4(KEYINPUT55), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n612_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(KEYINPUT56), .A3(new_n612_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n845_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n635_), .A2(new_n636_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n649_), .B1(new_n642_), .B2(new_n647_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859_));
  OR3_X1    g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n653_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n640_), .A2(new_n649_), .A3(new_n642_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n859_), .B1(new_n858_), .B2(new_n653_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n658_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n857_), .A2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n676_), .B1(new_n856_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n631_), .A2(new_n612_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n764_), .A2(new_n869_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n851_), .A2(KEYINPUT56), .A3(new_n612_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT56), .B1(new_n851_), .B2(new_n612_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n870_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n857_), .A2(new_n864_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT57), .A3(new_n676_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n864_), .A2(new_n869_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT58), .B(new_n877_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n716_), .A3(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n868_), .A2(new_n876_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n844_), .B1(new_n883_), .B2(new_n709_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n450_), .A2(new_n666_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n452_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n884_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G113gat), .B1(new_n889_), .B2(new_n662_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n880_), .A2(new_n716_), .A3(new_n881_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n875_), .B2(new_n676_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT118), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n868_), .A2(new_n894_), .A3(new_n882_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n893_), .A2(new_n876_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n844_), .B1(new_n896_), .B2(new_n709_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n888_), .A2(KEYINPUT59), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT59), .B1(new_n884_), .B2(new_n888_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n662_), .A2(G113gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT119), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n890_), .B1(new_n902_), .B2(new_n904_), .ZN(G1340gat));
  INV_X1    g704(.A(new_n899_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n638_), .B(new_n901_), .C1(new_n897_), .C2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G120gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n909_));
  AOI21_X1  g708(.A(G120gat), .B1(new_n638_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT120), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n909_), .B2(G120gat), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n889_), .B(new_n911_), .C1(new_n910_), .C2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n908_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT121), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n908_), .A2(new_n917_), .A3(new_n914_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1341gat));
  AOI21_X1  g718(.A(G127gat), .B1(new_n889_), .B2(new_n518_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n518_), .A2(G127gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n902_), .B2(new_n921_), .ZN(G1342gat));
  AND4_X1   g721(.A1(G134gat), .A2(new_n900_), .A3(new_n716_), .A4(new_n901_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G134gat), .B1(new_n889_), .B2(new_n593_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1343gat));
  NOR2_X1   g724(.A1(new_n884_), .A2(new_n453_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n885_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n662_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n638_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g731(.A1(new_n927_), .A2(new_n709_), .ZN(new_n933_));
  XOR2_X1   g732(.A(KEYINPUT61), .B(G155gat), .Z(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1346gat));
  AND3_X1   g734(.A1(new_n928_), .A2(G162gat), .A3(new_n716_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n927_), .A2(new_n676_), .ZN(new_n937_));
  OR3_X1    g736(.A1(new_n937_), .A2(KEYINPUT122), .A3(G162gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(KEYINPUT122), .B1(new_n937_), .B2(G162gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n936_), .B1(new_n938_), .B2(new_n939_), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n673_), .A2(new_n441_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n942_), .A2(new_n359_), .A3(new_n701_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n897_), .A2(new_n764_), .A3(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n291_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(KEYINPUT123), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n947_), .A2(KEYINPUT123), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n946_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n945_), .A2(new_n294_), .ZN(new_n951_));
  OAI211_X1 g750(.A(KEYINPUT123), .B(new_n947_), .C1(new_n945_), .C2(new_n291_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(G1348gat));
  NOR4_X1   g752(.A1(new_n884_), .A2(new_n607_), .A3(new_n639_), .A4(new_n944_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n897_), .A2(new_n944_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n638_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n956_), .B2(new_n290_), .ZN(G1349gat));
  INV_X1    g756(.A(new_n955_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n958_), .A2(new_n709_), .A3(new_n368_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n884_), .A2(new_n709_), .A3(new_n944_), .ZN(new_n960_));
  XOR2_X1   g759(.A(new_n960_), .B(KEYINPUT124), .Z(new_n961_));
  NOR2_X1   g760(.A1(new_n333_), .A2(new_n334_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n959_), .B1(new_n961_), .B2(new_n963_), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n958_), .B2(new_n715_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n955_), .A2(new_n367_), .A3(new_n593_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1351gat));
  NOR3_X1   g766(.A1(new_n884_), .A2(new_n453_), .A3(new_n942_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n662_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n638_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(KEYINPUT125), .B(G204gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1353gat));
  NAND2_X1  g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n968_), .A2(new_n518_), .A3(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(KEYINPUT126), .ZN(new_n976_));
  NOR2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978_));
  NAND4_X1  g777(.A1(new_n968_), .A2(new_n978_), .A3(new_n518_), .A4(new_n974_), .ZN(new_n979_));
  AND3_X1   g778(.A1(new_n976_), .A2(new_n977_), .A3(new_n979_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n977_), .B1(new_n976_), .B2(new_n979_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n980_), .A2(new_n981_), .ZN(G1354gat));
  NAND2_X1  g781(.A1(new_n968_), .A2(new_n716_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(KEYINPUT127), .B(G218gat), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n968_), .A2(new_n593_), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n985_), .B1(new_n986_), .B2(new_n984_), .ZN(G1355gat));
endmodule


