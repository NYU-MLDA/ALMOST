//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n982_,
    new_n983_, new_n984_;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n205_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT89), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n215_), .B(new_n216_), .C1(new_n209_), .C2(KEYINPUT2), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n202_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n223_));
  INV_X1    g022(.A(G197gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT92), .B1(new_n224_), .B2(G204gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT90), .B(G197gat), .Z(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(G204gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT90), .B(G197gat), .ZN(new_n228_));
  INV_X1    g027(.A(G204gat), .ZN(new_n229_));
  NOR3_X1   g028(.A1(new_n228_), .A2(KEYINPUT92), .A3(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n223_), .B1(new_n227_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT94), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(KEYINPUT94), .B(new_n223_), .C1(new_n227_), .C2(new_n230_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G211gat), .B(G218gat), .Z(new_n235_));
  OR3_X1    g034(.A1(new_n229_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT91), .B1(new_n229_), .B2(G197gat), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n236_), .B(new_n237_), .C1(new_n226_), .C2(G204gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n235_), .B1(new_n238_), .B2(KEYINPUT21), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n227_), .A2(new_n230_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(KEYINPUT21), .A3(new_n235_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n222_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n220_), .B(KEYINPUT28), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G228gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(G78gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G106gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G22gat), .B(G50gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n249_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n245_), .A2(new_n248_), .A3(new_n256_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261_));
  INV_X1    g060(.A(G120gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G113gat), .ZN(new_n263_));
  INV_X1    g062(.A(G113gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G120gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n265_), .A3(KEYINPUT87), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT87), .B1(new_n263_), .B2(new_n265_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n261_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT87), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n264_), .A2(G120gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n262_), .A2(G113gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n261_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n266_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT88), .B1(new_n269_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT88), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n267_), .A2(new_n268_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(new_n274_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n276_), .A2(new_n279_), .A3(KEYINPUT31), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G71gat), .B(G99gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT31), .B1(new_n276_), .B2(new_n279_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n284_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n286_), .B2(new_n280_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT86), .B(G43gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(G169gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(new_n293_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n292_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n293_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT84), .B1(new_n296_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n294_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n296_), .A2(KEYINPUT84), .A3(new_n300_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT25), .B(G183gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT81), .B1(new_n307_), .B2(G190gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT26), .B(G190gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n306_), .B(new_n308_), .C1(new_n309_), .C2(KEYINPUT81), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(G169gat), .B2(G176gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT82), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(G169gat), .B2(G176gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n314_), .A2(new_n316_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n310_), .B(new_n317_), .C1(KEYINPUT24), .C2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n299_), .B1(new_n305_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT85), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(KEYINPUT85), .B(new_n299_), .C1(new_n305_), .C2(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G227gat), .A2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(G15gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT30), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n327_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n290_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n322_), .A2(new_n323_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n327_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n290_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n328_), .A3(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n289_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n289_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n260_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n245_), .A2(new_n248_), .A3(new_n256_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n256_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n331_), .A2(new_n336_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n288_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n289_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT99), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n276_), .A2(new_n279_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT98), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .A4(new_n219_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n267_), .A2(new_n268_), .A3(new_n261_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n274_), .B1(new_n273_), .B2(new_n266_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n277_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n273_), .A2(new_n266_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT88), .B1(new_n356_), .B2(new_n261_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n355_), .A2(new_n357_), .A3(new_n219_), .A4(new_n351_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT98), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n352_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n355_), .A2(new_n219_), .A3(new_n357_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n211_), .B(new_n218_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(KEYINPUT4), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n348_), .B1(new_n360_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n364_), .A3(new_n362_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n352_), .A2(new_n359_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n369_), .A2(KEYINPUT99), .A3(new_n365_), .A4(new_n363_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G1gat), .B(G29gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G85gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT0), .B(G57gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n373_), .B(new_n374_), .Z(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n371_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n367_), .A2(new_n375_), .A3(new_n370_), .A4(new_n368_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n347_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n322_), .A2(new_n240_), .A3(new_n242_), .A4(new_n323_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT20), .ZN(new_n387_));
  INV_X1    g186(.A(new_n298_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n292_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT96), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT96), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(new_n392_), .A3(new_n292_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n297_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n309_), .A2(new_n306_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n317_), .A3(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n394_), .A2(new_n397_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n385_), .B1(new_n387_), .B2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G8gat), .B(G36gat), .Z(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT20), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n332_), .B2(new_n243_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n394_), .A2(new_n240_), .A3(new_n242_), .A4(new_n397_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n384_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n399_), .A2(new_n404_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT27), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n332_), .A2(new_n243_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n240_), .A2(new_n242_), .A3(new_n397_), .A4(new_n390_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(KEYINPUT20), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n385_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n393_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n392_), .B1(new_n389_), .B2(new_n292_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n397_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n243_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n418_), .A2(KEYINPUT20), .A3(new_n384_), .A4(new_n386_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n404_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT100), .B1(new_n410_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  INV_X1    g221(.A(new_n409_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n404_), .B1(new_n399_), .B2(new_n408_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n404_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n419_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n384_), .B1(new_n406_), .B2(new_n412_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT100), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT27), .A4(new_n409_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n421_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n381_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n337_), .A2(new_n338_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n342_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n423_), .A2(new_n424_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n378_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n378_), .A2(new_n438_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n369_), .A2(new_n364_), .A3(new_n363_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n361_), .A2(new_n365_), .A3(new_n362_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n376_), .A3(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n437_), .A2(new_n440_), .A3(new_n441_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n399_), .A2(new_n408_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n379_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n436_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n433_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G1gat), .B(G8gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT75), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455_));
  INV_X1    g254(.A(G1gat), .ZN(new_n456_));
  INV_X1    g255(.A(G8gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n453_), .A2(KEYINPUT75), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n453_), .A2(KEYINPUT75), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G29gat), .B(G36gat), .Z(new_n466_));
  XOR2_X1   g265(.A(G43gat), .B(G50gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT77), .B1(new_n465_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n454_), .A2(new_n459_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT77), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n468_), .A2(new_n471_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT76), .ZN(new_n480_));
  AOI211_X1 g279(.A(new_n480_), .B(new_n472_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT76), .B1(new_n476_), .B2(new_n478_), .ZN(new_n482_));
  OAI22_X1  g281(.A1(new_n473_), .A2(new_n479_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n481_), .A2(new_n482_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n478_), .B(KEYINPUT15), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n465_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n484_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n487_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n480_), .B1(new_n465_), .B2(new_n472_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n476_), .A2(KEYINPUT76), .A3(new_n478_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n485_), .B1(new_n489_), .B2(new_n465_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(KEYINPUT78), .A3(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n486_), .A2(new_n492_), .A3(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G113gat), .B(G141gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT79), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n486_), .A2(new_n492_), .A3(new_n497_), .A4(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT80), .Z(new_n507_));
  NOR2_X1   g306(.A1(new_n452_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G85gat), .B(G92gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OR3_X1    g310(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(G99gat), .B2(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n512_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT66), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n520_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT67), .B(new_n511_), .C1(new_n517_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT8), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n513_), .A2(G99gat), .A3(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n528_), .A2(new_n512_), .A3(new_n519_), .A4(new_n521_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n511_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT68), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n524_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n529_), .A2(KEYINPUT67), .A3(new_n511_), .A4(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n535_));
  INV_X1    g334(.A(G85gat), .ZN(new_n536_));
  OR2_X1    g335(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n535_), .B1(new_n539_), .B2(KEYINPUT9), .ZN(new_n540_));
  OR2_X1    g339(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(KEYINPUT64), .A3(new_n253_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n253_), .A3(new_n542_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT64), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n545_), .A2(new_n546_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n540_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n525_), .A2(new_n532_), .A3(new_n534_), .A4(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G71gat), .B(G78gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(KEYINPUT11), .ZN(new_n552_));
  INV_X1    g351(.A(new_n551_), .ZN(new_n553_));
  INV_X1    g352(.A(G64gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G57gat), .ZN(new_n555_));
  INV_X1    g354(.A(G57gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G64gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n557_), .A3(KEYINPUT11), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n552_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT69), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n563_), .B(new_n552_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n549_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n549_), .A2(new_n565_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n509_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n561_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n568_), .A2(new_n570_), .B1(new_n549_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n509_), .ZN(new_n574_));
  AND4_X1   g373(.A1(new_n525_), .A2(new_n532_), .A3(new_n534_), .A4(new_n548_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n565_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n569_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT5), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT70), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n578_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT13), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT35), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n549_), .A2(new_n489_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n590_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n549_), .B2(new_n472_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n591_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n575_), .A2(new_n478_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n591_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n549_), .A2(new_n489_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .A4(new_n593_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(KEYINPUT36), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n595_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT72), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n595_), .A2(new_n599_), .A3(KEYINPUT72), .A4(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n595_), .A2(new_n599_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n602_), .B(KEYINPUT36), .Z(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n608_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n606_), .A2(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n613_), .B(KEYINPUT74), .C1(new_n614_), .C2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT74), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n617_), .A3(new_n612_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n465_), .B(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(new_n561_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT17), .ZN(new_n623_));
  XOR2_X1   g422(.A(G127gat), .B(G155gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT16), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n622_), .A2(new_n623_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n561_), .B2(new_n621_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n627_), .B(new_n623_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n565_), .B2(new_n621_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(new_n565_), .B2(new_n621_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n586_), .A2(new_n619_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n508_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n456_), .A3(new_n379_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n506_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n586_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n399_), .A2(new_n408_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n426_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n441_), .A2(new_n643_), .A3(new_n409_), .A4(new_n444_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n450_), .B1(new_n644_), .B2(new_n439_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n436_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n379_), .B1(new_n339_), .B2(new_n346_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(new_n421_), .A3(new_n425_), .A4(new_n431_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n633_), .A2(new_n615_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n641_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n380_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n637_), .A2(new_n638_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n639_), .A2(new_n654_), .A3(new_n655_), .ZN(G1324gat));
  NAND3_X1  g455(.A1(new_n636_), .A2(new_n457_), .A3(new_n432_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n457_), .B1(new_n652_), .B2(new_n432_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n659_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n657_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT40), .B(new_n657_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1325gat));
  OAI21_X1  g468(.A(G15gat), .B1(new_n653_), .B2(new_n435_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n671_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n636_), .A2(new_n325_), .A3(new_n434_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(G1326gat));
  INV_X1    g474(.A(G22gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n652_), .B2(new_n260_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT42), .Z(new_n678_));
  NAND3_X1  g477(.A1(new_n636_), .A2(new_n676_), .A3(new_n260_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n633_), .A2(new_n615_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n586_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n508_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n379_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n619_), .A2(KEYINPUT103), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n687_), .A2(new_n689_), .B1(new_n433_), .B2(new_n451_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT43), .B1(new_n647_), .B2(new_n649_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n690_), .A2(KEYINPUT43), .B1(new_n691_), .B2(new_n619_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n641_), .A2(new_n633_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n686_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n693_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n619_), .B(KEYINPUT103), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n650_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n650_), .A2(new_n696_), .A3(new_n619_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n695_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n694_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n379_), .A2(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n685_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(new_n432_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n683_), .A2(G36gat), .A3(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT45), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n694_), .A2(new_n701_), .A3(new_n432_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n708_), .A2(KEYINPUT104), .A3(G36gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT104), .B1(new_n708_), .B2(G36gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n707_), .B(new_n712_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  NAND4_X1  g515(.A1(new_n694_), .A2(new_n701_), .A3(G43gat), .A4(new_n434_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n717_), .A2(KEYINPUT106), .ZN(new_n718_));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n683_), .B2(new_n435_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(KEYINPUT106), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT47), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n718_), .A2(new_n724_), .A3(new_n720_), .A4(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1330gat));
  AOI21_X1  g525(.A(G50gat), .B1(new_n684_), .B2(new_n260_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n260_), .A2(G50gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n702_), .B2(new_n728_), .ZN(G1331gat));
  NOR2_X1   g528(.A1(new_n452_), .A2(new_n506_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n633_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n619_), .ZN(new_n732_));
  AND4_X1   g531(.A1(new_n586_), .A2(new_n730_), .A3(new_n731_), .A4(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n556_), .A3(new_n379_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n650_), .A2(new_n507_), .A3(new_n586_), .A4(new_n651_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n380_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n735_), .B2(new_n705_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n432_), .A2(new_n554_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT107), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n733_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n735_), .B2(new_n435_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT49), .ZN(new_n745_));
  INV_X1    g544(.A(G71gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n733_), .A2(new_n746_), .A3(new_n434_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1334gat));
  OAI21_X1  g547(.A(G78gat), .B1(new_n735_), .B2(new_n342_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT50), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n733_), .A2(new_n251_), .A3(new_n260_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1335gat));
  NOR2_X1   g551(.A1(new_n585_), .A2(new_n681_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n730_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT108), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n536_), .A3(new_n379_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n692_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n586_), .A2(new_n640_), .A3(new_n633_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT109), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n379_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n756_), .B1(new_n761_), .B2(new_n536_), .ZN(G1336gat));
  AOI21_X1  g561(.A(G92gat), .B1(new_n755_), .B2(new_n432_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n705_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT110), .Z(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n760_), .B2(new_n765_), .ZN(G1337gat));
  NAND2_X1  g565(.A1(new_n760_), .A2(new_n434_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G99gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n755_), .A2(new_n434_), .A3(new_n543_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g570(.A1(new_n755_), .A2(new_n253_), .A3(new_n260_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n759_), .B(new_n260_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G106gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G106gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g577(.A1(new_n432_), .A2(new_n380_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n346_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n509_), .B1(new_n573_), .B2(new_n567_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n568_), .A2(new_n570_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n572_), .A2(new_n549_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n577_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT55), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n573_), .A2(new_n789_), .A3(new_n577_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n784_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n582_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n783_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n783_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT113), .B1(new_n791_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n785_), .A2(new_n786_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n574_), .B1(new_n797_), .B2(new_n566_), .ZN(new_n798_));
  AND4_X1   g597(.A1(new_n789_), .A2(new_n577_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n789_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n794_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n793_), .A2(new_n796_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n578_), .A2(new_n792_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n506_), .A2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n804_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n805_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n483_), .A2(new_n484_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n495_), .A2(new_n485_), .A3(new_n490_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n502_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n505_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT115), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n505_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n584_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n808_), .A2(new_n809_), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n782_), .B1(new_n820_), .B2(new_n615_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n804_), .A2(new_n807_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT114), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n804_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n818_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n615_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT116), .B1(new_n791_), .B2(new_n795_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n801_), .A2(new_n830_), .A3(new_n794_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n793_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n578_), .A2(new_n792_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n828_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n619_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n828_), .B(KEYINPUT58), .C1(new_n832_), .C2(new_n834_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT118), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n505_), .A2(new_n815_), .A3(new_n812_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n815_), .B1(new_n505_), .B2(new_n812_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n806_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT56), .B1(new_n801_), .B2(new_n582_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n830_), .B1(new_n801_), .B2(new_n794_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n845_), .B2(new_n831_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT58), .B1(new_n846_), .B2(new_n828_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n835_), .A2(new_n836_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n619_), .A4(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n821_), .A2(new_n827_), .A3(new_n839_), .A4(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT119), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n822_), .A2(KEYINPUT114), .B1(new_n584_), .B2(new_n817_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n782_), .B(new_n615_), .C1(new_n853_), .C2(new_n824_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT57), .B1(new_n825_), .B2(new_n826_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n839_), .A2(new_n850_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n852_), .A2(new_n859_), .A3(new_n633_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n861_));
  NAND4_X1  g660(.A1(new_n634_), .A2(KEYINPUT112), .A3(new_n507_), .A4(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n732_), .A2(new_n507_), .A3(new_n585_), .A4(new_n731_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n861_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n865_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n862_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n781_), .B1(new_n860_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n506_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n264_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n821_), .B(new_n827_), .C1(new_n838_), .C2(new_n837_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n633_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n868_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n872_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n507_), .A2(new_n264_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT120), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n877_), .B(new_n879_), .C1(new_n869_), .C2(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n871_), .A2(new_n881_), .ZN(G1340gat));
  OAI211_X1 g681(.A(new_n586_), .B(new_n877_), .C1(new_n869_), .C2(new_n880_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n262_), .B1(new_n585_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n869_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n262_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1341gat));
  OAI211_X1 g686(.A(new_n731_), .B(new_n877_), .C1(new_n869_), .C2(new_n880_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G127gat), .ZN(new_n889_));
  INV_X1    g688(.A(G127gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n869_), .A2(new_n890_), .A3(new_n731_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1342gat));
  OAI211_X1 g691(.A(new_n619_), .B(new_n877_), .C1(new_n869_), .C2(new_n880_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G134gat), .ZN(new_n894_));
  INV_X1    g693(.A(G134gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n869_), .A2(new_n895_), .A3(new_n615_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1343gat));
  AOI21_X1  g696(.A(new_n731_), .B1(new_n851_), .B2(KEYINPUT119), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n876_), .B1(new_n898_), .B2(new_n859_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n339_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n779_), .A2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT121), .B(G141gat), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n902_), .A2(new_n506_), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(new_n506_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1344gat));
  XNOR2_X1  g705(.A(KEYINPUT122), .B(G148gat), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n902_), .A2(new_n586_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n902_), .B2(new_n586_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1345gat));
  XNOR2_X1  g709(.A(KEYINPUT61), .B(G155gat), .ZN(new_n911_));
  INV_X1    g710(.A(new_n902_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n633_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n911_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n902_), .A2(new_n731_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1346gat));
  NAND2_X1  g715(.A1(new_n860_), .A2(new_n868_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n901_), .ZN(new_n918_));
  AND4_X1   g717(.A1(G162gat), .A2(new_n917_), .A3(new_n697_), .A4(new_n918_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n899_), .A2(new_n826_), .A3(new_n901_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT123), .B1(new_n920_), .B2(G162gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n917_), .A2(new_n615_), .A3(new_n918_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923_));
  INV_X1    g722(.A(G162gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n919_), .B1(new_n921_), .B2(new_n925_), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n705_), .A2(new_n379_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n346_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n874_), .B2(new_n868_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT22), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n931_), .A2(new_n932_), .A3(new_n506_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n933_), .A2(G169gat), .A3(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(G169gat), .ZN(new_n937_));
  INV_X1    g736(.A(new_n931_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n640_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n939_), .B2(new_n934_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n933_), .A2(new_n935_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n936_), .B1(new_n940_), .B2(new_n941_), .ZN(G1348gat));
  AOI21_X1  g741(.A(G176gat), .B1(new_n931_), .B2(new_n586_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n917_), .A2(new_n342_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n928_), .A2(new_n435_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n947_), .A2(G176gat), .A3(new_n586_), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n944_), .B(new_n945_), .C1(new_n946_), .C2(new_n948_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n899_), .A2(new_n260_), .A3(new_n948_), .ZN(new_n950_));
  OAI21_X1  g749(.A(KEYINPUT125), .B1(new_n950_), .B2(new_n943_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n951_), .ZN(G1349gat));
  NOR3_X1   g751(.A1(new_n938_), .A2(new_n306_), .A3(new_n633_), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n917_), .A2(new_n342_), .A3(new_n731_), .A4(new_n947_), .ZN(new_n954_));
  INV_X1    g753(.A(G183gat), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n953_), .B1(new_n954_), .B2(new_n955_), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n938_), .B2(new_n732_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n931_), .A2(new_n309_), .A3(new_n615_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n928_), .A2(new_n339_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n917_), .A2(new_n960_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n961_), .A2(new_n224_), .A3(new_n640_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n960_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n899_), .A2(new_n963_), .ZN(new_n964_));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964_), .B2(new_n506_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n962_), .A2(new_n965_), .ZN(G1352gat));
  OAI21_X1  g765(.A(G204gat), .B1(new_n961_), .B2(new_n585_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n964_), .A2(new_n229_), .A3(new_n586_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(G1353gat));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n970_));
  INV_X1    g769(.A(G211gat), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n970_), .A2(new_n971_), .A3(KEYINPUT126), .ZN(new_n972_));
  XOR2_X1   g771(.A(new_n972_), .B(KEYINPUT127), .Z(new_n973_));
  INV_X1    g772(.A(new_n973_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n731_), .B1(new_n970_), .B2(new_n971_), .ZN(new_n975_));
  NOR3_X1   g774(.A1(new_n899_), .A2(new_n963_), .A3(new_n975_), .ZN(new_n976_));
  AOI21_X1  g775(.A(KEYINPUT126), .B1(new_n970_), .B2(new_n971_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n974_), .B1(new_n976_), .B2(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n977_), .ZN(new_n979_));
  OAI211_X1 g778(.A(new_n979_), .B(new_n973_), .C1(new_n961_), .C2(new_n975_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n978_), .A2(new_n980_), .ZN(G1354gat));
  OAI21_X1  g780(.A(G218gat), .B1(new_n961_), .B2(new_n732_), .ZN(new_n982_));
  INV_X1    g781(.A(G218gat), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n964_), .A2(new_n983_), .A3(new_n615_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n982_), .A2(new_n984_), .ZN(G1355gat));
endmodule


