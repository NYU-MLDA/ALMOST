//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT83), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT85), .Z(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT3), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT86), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(KEYINPUT1), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n217_), .A2(KEYINPUT84), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n217_), .B(KEYINPUT84), .C1(KEYINPUT1), .C2(new_n215_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n209_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n204_), .A4(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n202_), .B1(new_n214_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G211gat), .B(G218gat), .Z(new_n224_));
  INV_X1    g023(.A(G197gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G204gat), .ZN(new_n226_));
  INV_X1    g025(.A(G204gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G197gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n224_), .A2(KEYINPUT21), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT89), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(new_n224_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n226_), .A2(new_n228_), .A3(KEYINPUT88), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n234_), .B(KEYINPUT21), .C1(KEYINPUT88), .C2(new_n226_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(G228gat), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n223_), .A2(new_n237_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n241_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n237_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(new_n222_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G78gat), .B(G106gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n214_), .A2(new_n221_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(KEYINPUT29), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G22gat), .B(G50gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT28), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n252_), .B(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n242_), .A2(new_n245_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n246_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n248_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n258_), .A2(KEYINPUT90), .A3(new_n248_), .A4(new_n255_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT19), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT24), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  MUX2_X1   g066(.A(new_n266_), .B(KEYINPUT24), .S(new_n267_), .Z(new_n268_));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT23), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT25), .B(G183gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(new_n272_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n244_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n269_), .A2(new_n270_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n265_), .B(KEYINPUT93), .Z(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT81), .B(G176gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT22), .B(G169gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT94), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n282_), .A2(KEYINPUT94), .A3(new_n285_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n281_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n277_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT78), .B(G190gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(G183gat), .ZN(new_n293_));
  INV_X1    g092(.A(G169gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT22), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT79), .ZN(new_n296_));
  OR3_X1    g095(.A1(new_n294_), .A2(KEYINPUT80), .A3(KEYINPUT22), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT80), .B1(new_n294_), .B2(KEYINPUT22), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n283_), .A3(new_n298_), .ZN(new_n299_));
  OAI221_X1 g098(.A(new_n265_), .B1(new_n293_), .B2(new_n271_), .C1(new_n296_), .C2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n273_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n292_), .B2(KEYINPUT26), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n268_), .B(new_n272_), .C1(new_n301_), .C2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n237_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n264_), .B1(new_n291_), .B2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n231_), .A2(new_n300_), .A3(new_n236_), .A4(new_n304_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT91), .B1(new_n310_), .B2(KEYINPUT20), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT92), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n276_), .A2(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n268_), .A2(new_n272_), .A3(KEYINPUT92), .A4(new_n275_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(new_n290_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n312_), .B(new_n313_), .C1(new_n318_), .C2(new_n244_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n309_), .B1(new_n319_), .B2(new_n264_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT18), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n313_), .B1(new_n244_), .B2(new_n318_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n264_), .B1(new_n327_), .B2(new_n311_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n318_), .A2(new_n244_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT20), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n264_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n306_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n324_), .A3(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n326_), .A2(KEYINPUT27), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT102), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT102), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n326_), .A2(new_n336_), .A3(KEYINPUT27), .A4(new_n333_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT95), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n333_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n328_), .A2(new_n332_), .A3(KEYINPUT95), .A4(new_n324_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n328_), .A2(new_n332_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n325_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT27), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G1gat), .B(G29gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G57gat), .B(G85gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G127gat), .B(G134gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT82), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n353_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n355_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT4), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n251_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT97), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n251_), .A2(new_n361_), .A3(KEYINPUT97), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n352_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n356_), .A2(new_n360_), .ZN(new_n367_));
  OR3_X1    g166(.A1(new_n251_), .A2(KEYINPUT96), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n251_), .B2(KEYINPUT96), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(KEYINPUT4), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT98), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n369_), .A3(new_n352_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n351_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n351_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n373_), .A4(new_n372_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G43gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n305_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(new_n367_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(G15gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT30), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT31), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n384_), .B(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n380_), .A2(new_n390_), .ZN(new_n391_));
  AND4_X1   g190(.A1(new_n262_), .A2(new_n338_), .A3(new_n346_), .A4(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n390_), .ZN(new_n393_));
  AND4_X1   g192(.A1(new_n376_), .A2(new_n379_), .A3(new_n261_), .A4(new_n260_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n394_), .A2(new_n346_), .A3(new_n335_), .A4(new_n337_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n393_), .B1(new_n396_), .B2(KEYINPUT103), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT103), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n379_), .A2(KEYINPUT33), .ZN(new_n399_));
  INV_X1    g198(.A(new_n374_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n378_), .A4(new_n377_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n352_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n368_), .A2(new_n369_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n351_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT100), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT100), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n408_), .A3(new_n351_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n404_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n370_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n412_));
  AND4_X1   g211(.A1(new_n341_), .A2(new_n340_), .A3(new_n343_), .A4(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n324_), .A2(KEYINPUT32), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n342_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n320_), .B2(new_n414_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n403_), .A2(new_n413_), .B1(new_n380_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n262_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n395_), .B(new_n398_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n392_), .B1(new_n397_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G120gat), .B(G148gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT5), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G176gat), .B(G204gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n422_), .B(new_n423_), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT66), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT64), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT6), .ZN(new_n430_));
  AND2_X1   g229(.A1(G99gat), .A2(G106gat), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n434_));
  INV_X1    g233(.A(G99gat), .ZN(new_n435_));
  INV_X1    g234(.A(G106gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n432_), .A2(new_n433_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G85gat), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n426_), .B1(new_n440_), .B2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n429_), .A2(KEYINPUT6), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n427_), .A2(KEYINPUT64), .ZN(new_n448_));
  OAI22_X1  g247(.A1(new_n447_), .A2(new_n448_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n437_), .A2(new_n438_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n445_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(KEYINPUT66), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(KEYINPUT8), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n426_), .B(new_n456_), .C1(new_n440_), .C2(new_n445_), .ZN(new_n457_));
  OR2_X1    g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n436_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n443_), .A2(KEYINPUT9), .A3(new_n444_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n444_), .A2(KEYINPUT9), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n432_), .A2(new_n433_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT65), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT65), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n449_), .A2(new_n451_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n455_), .A2(new_n457_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G64gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G57gat), .ZN(new_n473_));
  INV_X1    g272(.A(G57gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G64gat), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G71gat), .B(G78gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(KEYINPUT11), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n476_), .A2(KEYINPUT11), .ZN(new_n479_));
  INV_X1    g278(.A(new_n477_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n473_), .A2(new_n475_), .A3(KEYINPUT11), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n478_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT12), .B1(new_n471_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G230gat), .A2(G233gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n455_), .A2(new_n470_), .A3(new_n457_), .A4(new_n483_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n483_), .A2(KEYINPUT67), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(new_n478_), .C1(new_n479_), .C2(new_n482_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n489_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n446_), .A2(KEYINPUT8), .A3(new_n454_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n457_), .A2(new_n469_), .A3(new_n465_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .A4(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n487_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n488_), .ZN(new_n499_));
  AOI211_X1 g298(.A(KEYINPUT66), .B(KEYINPUT8), .C1(new_n452_), .C2(new_n453_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n465_), .A2(new_n469_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n483_), .B1(new_n502_), .B2(new_n455_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n499_), .B2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n425_), .B1(new_n497_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n488_), .B(new_n496_), .C1(new_n503_), .C2(KEYINPUT12), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n504_), .B(new_n425_), .C1(new_n507_), .C2(new_n498_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT69), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n506_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n509_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT69), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n505_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT13), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(new_n517_), .A3(KEYINPUT13), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT70), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n524_), .A3(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n527_));
  XOR2_X1   g326(.A(G29gat), .B(G36gat), .Z(new_n528_));
  XOR2_X1   g327(.A(G43gat), .B(G50gat), .Z(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G29gat), .B(G36gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G43gat), .B(G50gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT75), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(KEYINPUT75), .A3(new_n533_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539_));
  INV_X1    g338(.A(G1gat), .ZN(new_n540_));
  INV_X1    g339(.A(G8gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT14), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G1gat), .B(G8gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT72), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(KEYINPUT72), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n543_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n543_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n545_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n538_), .A2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n536_), .A2(new_n551_), .A3(new_n537_), .A4(new_n548_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(KEYINPUT76), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n538_), .A2(new_n558_), .A3(new_n552_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n534_), .B(KEYINPUT15), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n552_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(new_n556_), .A3(new_n554_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G169gat), .B(G197gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n527_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(KEYINPUT77), .A3(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n420_), .A2(new_n526_), .A3(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n471_), .A2(new_n561_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT34), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n534_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n471_), .B2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT71), .B(new_n580_), .C1(new_n471_), .C2(new_n581_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n578_), .A2(new_n579_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n584_), .B(new_n585_), .C1(new_n575_), .C2(new_n582_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(KEYINPUT36), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n589_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n592_), .B(KEYINPUT36), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT37), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n589_), .A2(new_n596_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n600_), .B(new_n601_), .C1(new_n594_), .C2(new_n589_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT17), .ZN(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n552_), .B(new_n610_), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT73), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n490_), .A2(new_n492_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n604_), .B(new_n609_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n614_), .B1(new_n613_), .B2(new_n612_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n611_), .A2(new_n483_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n611_), .A2(new_n483_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n609_), .B(KEYINPUT17), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n603_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n574_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n540_), .A3(new_n380_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT38), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n526_), .A2(new_n573_), .A3(new_n620_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n625_), .A2(KEYINPUT104), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n595_), .A2(new_n598_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n420_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(KEYINPUT104), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n626_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n630_), .A2(new_n380_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n624_), .B1(new_n540_), .B2(new_n631_), .ZN(G1324gat));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n338_), .A2(new_n346_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n626_), .A2(new_n634_), .A3(new_n628_), .A4(new_n629_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n634_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(G8gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n574_), .A2(new_n621_), .A3(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT105), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT39), .B1(new_n635_), .B2(G8gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n633_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n644_), .A2(KEYINPUT40), .A3(new_n636_), .A4(new_n640_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1325gat));
  NAND3_X1  g445(.A1(new_n622_), .A2(new_n386_), .A3(new_n393_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n630_), .A2(new_n393_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n648_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT41), .B1(new_n648_), .B2(G15gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n622_), .A2(new_n652_), .A3(new_n418_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n630_), .A2(new_n418_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(G22gat), .ZN(new_n656_));
  AOI211_X1 g455(.A(KEYINPUT42), .B(new_n652_), .C1(new_n630_), .C2(new_n418_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(G1327gat));
  INV_X1    g457(.A(new_n620_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n627_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n380_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(G29gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n574_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n599_), .A2(new_n602_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n665_), .B2(KEYINPUT106), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n420_), .B2(new_n665_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n338_), .A2(new_n262_), .A3(new_n346_), .A4(new_n391_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n395_), .A2(new_n398_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n403_), .A2(new_n413_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n416_), .A2(new_n380_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n418_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n390_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n669_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n603_), .A3(new_n666_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n668_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n573_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n523_), .A2(new_n679_), .A3(new_n525_), .A4(new_n620_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n678_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n683_), .B(new_n680_), .C1(new_n668_), .C2(new_n677_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n380_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G29gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n685_), .B2(new_n380_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n664_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n685_), .B2(new_n634_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n574_), .A2(new_n692_), .A3(new_n634_), .A4(new_n661_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT45), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n682_), .A2(new_n684_), .A3(new_n637_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n695_), .B(KEYINPUT46), .C1(new_n698_), .C2(new_n692_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1329gat));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(G43gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n685_), .B2(new_n393_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n574_), .A2(new_n702_), .A3(new_n393_), .A4(new_n661_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n682_), .A2(new_n684_), .A3(new_n390_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT47), .B(new_n704_), .C1(new_n707_), .C2(new_n702_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1330gat));
  INV_X1    g508(.A(G50gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n262_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n574_), .A2(new_n418_), .A3(new_n661_), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n685_), .A2(new_n711_), .B1(new_n712_), .B2(new_n710_), .ZN(G1331gat));
  NOR2_X1   g512(.A1(new_n420_), .A2(new_n679_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(new_n526_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n621_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n380_), .A3(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n679_), .B(new_n620_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n628_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT109), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n662_), .A2(new_n474_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n719_), .A2(new_n474_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  NAND3_X1  g523(.A1(new_n716_), .A2(new_n472_), .A3(new_n634_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n722_), .A2(new_n634_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G64gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT48), .B(new_n472_), .C1(new_n722_), .C2(new_n634_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n716_), .A2(new_n731_), .A3(new_n393_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n722_), .A2(new_n393_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G71gat), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT49), .B(new_n731_), .C1(new_n722_), .C2(new_n393_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1334gat));
  INV_X1    g536(.A(G78gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n716_), .A2(new_n738_), .A3(new_n418_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n722_), .A2(new_n418_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G78gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT50), .B(new_n738_), .C1(new_n722_), .C2(new_n418_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1335gat));
  AND2_X1   g543(.A1(new_n715_), .A2(new_n661_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n441_), .A3(new_n380_), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n679_), .B(new_n659_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n678_), .A2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(new_n380_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(new_n441_), .ZN(G1336gat));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n442_), .A3(new_n634_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n748_), .A2(new_n634_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n442_), .ZN(G1337gat));
  NAND2_X1  g552(.A1(new_n748_), .A2(new_n393_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G99gat), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n745_), .A2(new_n458_), .A3(new_n459_), .A4(new_n393_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT51), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n756_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1338gat));
  NOR2_X1   g560(.A1(new_n262_), .A2(G106gat), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n714_), .A2(new_n526_), .A3(new_n661_), .A4(new_n762_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT110), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n678_), .A2(new_n418_), .A3(new_n747_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G106gat), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n764_), .A2(new_n768_), .A3(new_n772_), .A4(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  NOR2_X1   g573(.A1(new_n634_), .A2(new_n418_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n380_), .A3(new_n393_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT116), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n775_), .A2(new_n778_), .A3(new_n380_), .A4(new_n393_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n496_), .A2(new_n488_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(new_n485_), .A3(new_n498_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n498_), .B1(new_n781_), .B2(new_n485_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(KEYINPUT55), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n507_), .A2(new_n785_), .A3(new_n498_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n424_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT111), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n789_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n424_), .B(new_n791_), .C1(new_n784_), .C2(new_n786_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n570_), .A2(new_n572_), .A3(new_n508_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n790_), .A2(KEYINPUT112), .A3(new_n792_), .A4(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n554_), .A2(new_n557_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n566_), .B1(new_n796_), .B2(new_n562_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n555_), .A2(new_n556_), .A3(new_n559_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n567_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT113), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n567_), .A2(new_n799_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n513_), .A2(new_n517_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n795_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n793_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT112), .B1(new_n807_), .B2(new_n792_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n660_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT57), .B(new_n660_), .C1(new_n806_), .C2(new_n808_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT114), .B(KEYINPUT58), .Z(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n803_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n802_), .B1(new_n567_), .B2(new_n799_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n508_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n787_), .B2(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n783_), .A2(KEYINPUT55), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n497_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n786_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n425_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n788_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n815_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n813_), .B1(new_n825_), .B2(new_n665_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n824_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n497_), .A2(new_n504_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n828_), .A2(new_n425_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n823_), .B2(new_n788_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n787_), .A2(KEYINPUT56), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n814_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT115), .A3(new_n603_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n826_), .A2(new_n827_), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n811_), .A2(new_n812_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n620_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n603_), .A2(new_n679_), .A3(new_n620_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n837_), .A2(new_n522_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n837_), .B2(new_n522_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n780_), .B1(new_n836_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT117), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n841_), .B1(new_n620_), .B2(new_n835_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n846_), .B(KEYINPUT59), .C1(new_n847_), .C2(new_n780_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n836_), .A2(KEYINPUT118), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n835_), .A2(new_n851_), .A3(new_n620_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n841_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n780_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n844_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT119), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n835_), .A2(new_n851_), .A3(new_n620_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n851_), .B1(new_n835_), .B2(new_n620_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n842_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n844_), .A4(new_n854_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n849_), .A2(new_n856_), .A3(new_n679_), .A4(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G113gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n843_), .ZN(new_n864_));
  OR3_X1    g663(.A1(new_n864_), .A2(G113gat), .A3(new_n573_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1340gat));
  NAND4_X1  g665(.A1(new_n849_), .A2(new_n856_), .A3(new_n526_), .A4(new_n861_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G120gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT60), .B1(new_n523_), .B2(new_n525_), .ZN(new_n869_));
  MUX2_X1   g668(.A(new_n869_), .B(KEYINPUT60), .S(G120gat), .Z(new_n870_));
  NAND2_X1  g669(.A1(new_n843_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n620_), .A2(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT120), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n849_), .A2(new_n856_), .A3(new_n861_), .A4(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n873_), .B1(new_n864_), .B2(new_n620_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1342gat));
  NAND4_X1  g677(.A1(new_n849_), .A2(new_n856_), .A3(new_n603_), .A4(new_n861_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G134gat), .ZN(new_n880_));
  OR3_X1    g679(.A1(new_n864_), .A2(G134gat), .A3(new_n660_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n418_), .A2(new_n390_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n847_), .A2(new_n662_), .A3(new_n634_), .A4(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n679_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n526_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT121), .B(G148gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n884_), .A2(new_n659_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n884_), .B2(new_n627_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n603_), .A2(G162gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT122), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n884_), .B2(new_n895_), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n634_), .A2(new_n391_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n262_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n853_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n679_), .A2(new_n284_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT124), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n859_), .A2(new_n679_), .A3(new_n262_), .A4(new_n898_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  AND4_X1   g704(.A1(KEYINPUT123), .A2(new_n904_), .A3(new_n905_), .A4(G169gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n294_), .B1(new_n907_), .B2(KEYINPUT62), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n904_), .A2(new_n908_), .B1(KEYINPUT123), .B2(new_n905_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n903_), .B1(new_n906_), .B2(new_n909_), .ZN(G1348gat));
  NOR2_X1   g709(.A1(new_n847_), .A2(new_n418_), .ZN(new_n911_));
  AND4_X1   g710(.A1(G176gat), .A2(new_n911_), .A3(new_n526_), .A4(new_n898_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n900_), .A2(new_n526_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n283_), .ZN(G1349gat));
  NAND2_X1  g713(.A1(new_n898_), .A2(new_n659_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G183gat), .B1(new_n911_), .B2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n620_), .A2(new_n273_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n900_), .B2(new_n918_), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n900_), .A2(new_n274_), .A3(new_n627_), .ZN(new_n920_));
  INV_X1    g719(.A(G190gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n853_), .A2(new_n665_), .A3(new_n899_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1351gat));
  NAND2_X1  g722(.A1(new_n836_), .A2(new_n842_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n637_), .A2(new_n380_), .A3(new_n883_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI22_X1  g726(.A1(new_n927_), .A2(new_n573_), .B1(KEYINPUT125), .B2(new_n225_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n225_), .A2(KEYINPUT125), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT126), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n928_), .B(new_n930_), .ZN(G1352gat));
  NAND2_X1  g730(.A1(new_n926_), .A2(new_n526_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g732(.A(new_n620_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n926_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT127), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n926_), .A2(new_n938_), .A3(new_n934_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n936_), .A2(new_n937_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n937_), .B1(new_n936_), .B2(new_n939_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1354gat));
  OR3_X1    g741(.A1(new_n927_), .A2(G218gat), .A3(new_n660_), .ZN(new_n943_));
  OAI21_X1  g742(.A(G218gat), .B1(new_n927_), .B2(new_n665_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1355gat));
endmodule


