//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT64), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n207_), .A2(KEYINPUT65), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G85gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n208_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n206_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT10), .B(G99gat), .Z(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n220_), .A2(new_n221_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n219_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n209_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n223_), .A2(new_n225_), .ZN(new_n237_));
  AOI211_X1 g036(.A(new_n229_), .B(new_n232_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT7), .ZN(new_n239_));
  INV_X1    g038(.A(G99gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n221_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n224_), .B1(G99gat), .B2(G106gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n233_), .B(new_n241_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n209_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n228_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n227_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G29gat), .B(G36gat), .Z(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT70), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G29gat), .B(G36gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G43gat), .B(G50gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n204_), .B(new_n205_), .C1(new_n247_), .C2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT15), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n249_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n254_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n256_), .A2(KEYINPUT15), .A3(new_n257_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n247_), .A2(KEYINPUT68), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n227_), .B(new_n268_), .C1(new_n238_), .C2(new_n246_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n260_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n260_), .A2(new_n270_), .A3(KEYINPUT74), .ZN(new_n274_));
  INV_X1    g073(.A(new_n204_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n205_), .B1(new_n247_), .B2(new_n258_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(KEYINPUT71), .B(new_n205_), .C1(new_n247_), .C2(new_n258_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n270_), .A3(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n273_), .A2(new_n274_), .B1(new_n275_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G190gat), .B(G218gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT72), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G134gat), .B(G162gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT36), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT75), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n280_), .A2(new_n275_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n274_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT74), .B1(new_n260_), .B2(new_n270_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292_));
  INV_X1    g091(.A(new_n286_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT37), .ZN(new_n296_));
  INV_X1    g095(.A(new_n285_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n298_));
  AND2_X1   g097(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n291_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n295_), .A2(new_n296_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT76), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n287_), .B2(new_n294_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(KEYINPUT76), .A3(new_n296_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n302_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n305_), .A2(new_n307_), .B1(KEYINPUT37), .B2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G1gat), .B(G8gat), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G1gat), .A2(G8gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT14), .ZN(new_n313_));
  INV_X1    g112(.A(G15gat), .ZN(new_n314_));
  INV_X1    g113(.A(G22gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G15gat), .A2(G22gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n313_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(KEYINPUT77), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(KEYINPUT77), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n311_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(new_n310_), .A3(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(G71gat), .A2(G78gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G71gat), .A2(G78gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G57gat), .B(G64gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n332_), .B1(new_n333_), .B2(KEYINPUT11), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n333_), .B2(KEYINPUT11), .ZN(new_n336_));
  INV_X1    g135(.A(G64gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G57gat), .ZN(new_n338_));
  INV_X1    g137(.A(G57gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G64gat), .ZN(new_n340_));
  AND4_X1   g139(.A1(new_n335_), .A2(new_n338_), .A3(new_n340_), .A4(KEYINPUT11), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n334_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(new_n340_), .A3(KEYINPUT11), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT67), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(new_n340_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT11), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n338_), .A2(new_n340_), .A3(new_n335_), .A4(KEYINPUT11), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n344_), .A2(new_n347_), .A3(new_n332_), .A4(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n342_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G231gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n329_), .B(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G127gat), .B(G155gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G183gat), .B(G211gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT17), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(KEYINPUT17), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n353_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n353_), .A2(new_n359_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n309_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT80), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT83), .B(G169gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(G183gat), .B2(G190gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n369_), .A2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n371_), .A2(KEYINPUT82), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n371_), .A2(KEYINPUT82), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n373_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT25), .B(G183gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT26), .B(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(KEYINPUT24), .A3(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n384_), .A2(KEYINPUT24), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n380_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n390_), .B(G43gat), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n377_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  OAI22_X1  g192(.A1(new_n376_), .A2(new_n369_), .B1(new_n380_), .B2(new_n388_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n391_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(G15gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT30), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n396_), .B(new_n314_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT31), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n398_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n402_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n393_), .A2(new_n395_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT84), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT84), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n406_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G127gat), .B(G134gat), .Z(new_n413_));
  XOR2_X1   g212(.A(G113gat), .B(G120gat), .Z(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  AND3_X1   g214(.A1(new_n409_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT27), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G197gat), .B(G204gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT21), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G211gat), .B(G218gat), .Z(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n420_), .B(KEYINPUT21), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(new_n423_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n377_), .A2(new_n389_), .A3(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT22), .B(G169gat), .ZN(new_n428_));
  INV_X1    g227(.A(G176gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n385_), .B(new_n430_), .C1(new_n380_), .C2(new_n375_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n388_), .A2(new_n374_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT20), .B(new_n427_), .C1(new_n433_), .C2(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT19), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G8gat), .B(G36gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT18), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n431_), .A2(new_n432_), .A3(new_n426_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n431_), .A2(new_n432_), .A3(new_n426_), .A4(KEYINPUT92), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n436_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n448_), .A2(KEYINPUT20), .ZN(new_n449_));
  INV_X1    g248(.A(new_n424_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n420_), .A2(new_n421_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n423_), .B1(new_n422_), .B2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n453_), .A2(new_n394_), .A3(KEYINPUT91), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT91), .B1(new_n453_), .B2(new_n394_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n449_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n437_), .B(new_n441_), .C1(new_n447_), .C2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n455_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n394_), .A3(KEYINPUT91), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n441_), .B1(new_n462_), .B2(new_n437_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n419_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n434_), .A2(new_n436_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n442_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n448_), .B1(new_n461_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n465_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n454_), .A2(new_n455_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n436_), .B1(new_n472_), .B2(new_n467_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT94), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n441_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n457_), .A2(KEYINPUT27), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n418_), .B(new_n464_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G22gat), .B(G50gat), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G155gat), .B(G162gat), .Z(new_n480_));
  INV_X1    g279(.A(KEYINPUT1), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n483_));
  INV_X1    g282(.A(G141gat), .ZN(new_n484_));
  INV_X1    g283(.A(G148gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n485_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n482_), .A2(new_n483_), .A3(new_n487_), .A4(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n493_), .B(new_n495_), .C1(new_n486_), .C2(KEYINPUT2), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n480_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n489_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT28), .B1(new_n498_), .B2(KEYINPUT29), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT28), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT29), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n489_), .A2(new_n497_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n499_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n499_), .B2(new_n503_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n479_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n499_), .A2(new_n503_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT87), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n499_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n478_), .A3(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n510_), .A3(KEYINPUT90), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G78gat), .B(G106gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT89), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n513_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n506_), .A2(new_n510_), .A3(KEYINPUT90), .A4(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n506_), .A2(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n426_), .B1(KEYINPUT29), .B2(new_n498_), .ZN(new_n521_));
  AND2_X1   g320(.A1(G228gat), .A2(G233gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT88), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n521_), .B(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(KEYINPUT88), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n520_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n517_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n527_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G29gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G85gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT0), .B(G57gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(G225gat), .A2(G233gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n498_), .A2(new_n415_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n413_), .B(new_n414_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n489_), .A3(new_n497_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(KEYINPUT4), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT4), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n498_), .A2(new_n415_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n538_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n538_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n537_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n545_), .A2(new_n537_), .A3(new_n547_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n477_), .A2(new_n533_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n441_), .ZN(new_n554_));
  OAI22_X1  g353(.A1(new_n473_), .A2(KEYINPUT94), .B1(new_n436_), .B2(new_n434_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n469_), .A2(new_n470_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n476_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n437_), .B1(new_n447_), .B2(new_n456_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n554_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n457_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n557_), .A2(new_n558_), .B1(new_n561_), .B2(new_n419_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n533_), .A2(new_n562_), .A3(new_n551_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n441_), .A2(KEYINPUT32), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  OAI22_X1  g365(.A1(new_n549_), .A2(new_n550_), .B1(new_n559_), .B2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n542_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n537_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n539_), .A2(new_n546_), .A3(new_n541_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n560_), .A2(new_n571_), .A3(new_n457_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n548_), .B(new_n573_), .ZN(new_n574_));
  OAI22_X1  g373(.A1(new_n565_), .A2(new_n567_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n532_), .A3(new_n530_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n563_), .A2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n418_), .A2(KEYINPUT85), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n418_), .A2(KEYINPUT85), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n553_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n342_), .A2(new_n349_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n267_), .A2(new_n269_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n223_), .A2(new_n225_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n241_), .A2(new_n233_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n245_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n229_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n244_), .A2(new_n228_), .A3(new_n245_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n590_), .A2(new_n591_), .B1(new_n219_), .B2(new_n226_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n582_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n583_), .B1(new_n592_), .B2(new_n582_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n585_), .A2(new_n586_), .A3(new_n593_), .A4(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n586_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n247_), .A2(new_n350_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n590_), .A2(new_n591_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n582_), .B1(new_n598_), .B2(new_n227_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n595_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT5), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G176gat), .B(G204gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT69), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n601_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT13), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n258_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n326_), .A2(new_n328_), .A3(new_n266_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n326_), .A2(new_n328_), .A3(new_n258_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n617_), .B1(new_n615_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT81), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n619_), .A2(new_n621_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n617_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n620_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n614_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n626_), .B1(new_n618_), .B2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n613_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n581_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n366_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(G1gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n552_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n640_));
  XOR2_X1   g439(.A(new_n639_), .B(new_n640_), .Z(new_n641_));
  NOR2_X1   g440(.A1(new_n306_), .A2(new_n364_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT96), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n638_), .B1(new_n644_), .B2(new_n552_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n641_), .A2(new_n645_), .ZN(G1324gat));
  OAI21_X1  g445(.A(G8gat), .B1(new_n643_), .B2(new_n562_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT97), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT97), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(KEYINPUT39), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n647_), .A2(KEYINPUT97), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(G8gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n562_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n637_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n650_), .A2(new_n652_), .A3(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g456(.A(new_n580_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n314_), .B1(new_n644_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT41), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(KEYINPUT41), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n637_), .A2(new_n314_), .A3(new_n658_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(G1326gat));
  AOI21_X1  g463(.A(new_n315_), .B1(new_n644_), .B2(new_n533_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT42), .Z(new_n666_));
  NAND2_X1  g465(.A1(new_n533_), .A2(new_n315_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT98), .Z(new_n668_));
  NAND2_X1  g467(.A1(new_n637_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(new_n306_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n363_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n636_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(G29gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n676_), .A3(new_n552_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n635_), .A2(new_n363_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n308_), .A2(KEYINPUT37), .ZN(new_n680_));
  INV_X1    g479(.A(new_n307_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT76), .B1(new_n306_), .B2(new_n296_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n581_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n679_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n477_), .A2(new_n533_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n551_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n552_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n531_), .A2(new_n516_), .A3(new_n514_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n531_), .B1(new_n516_), .B2(new_n514_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n689_), .A2(new_n562_), .B1(new_n692_), .B2(new_n575_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n693_), .B2(new_n658_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n694_), .A2(new_n679_), .A3(new_n685_), .A4(new_n309_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n581_), .B2(new_n683_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n678_), .B1(new_n686_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n678_), .C1(new_n686_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n551_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT100), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G29gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n703_), .A2(KEYINPUT100), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n677_), .B1(new_n705_), .B2(new_n706_), .ZN(G1328gat));
  NOR2_X1   g506(.A1(new_n562_), .A2(G36gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n675_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT45), .ZN(new_n710_));
  INV_X1    g509(.A(G36gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n702_), .A2(new_n562_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n710_), .B(KEYINPUT46), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND2_X1  g516(.A1(new_n418_), .A2(G43gat), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n675_), .A2(new_n658_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT102), .B(G43gat), .Z(new_n720_));
  OAI22_X1  g519(.A1(new_n702_), .A2(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n675_), .A2(new_n723_), .A3(new_n533_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n700_), .A2(new_n533_), .A3(new_n701_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n725_), .A2(KEYINPUT103), .A3(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT103), .B1(new_n725_), .B2(G50gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT104), .B(new_n724_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n581_), .A2(new_n634_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n734_), .A2(KEYINPUT105), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n613_), .B1(new_n734_), .B2(KEYINPUT105), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n366_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n339_), .A3(new_n552_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n612_), .A3(new_n642_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n551_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1332gat));
  NAND3_X1  g541(.A1(new_n738_), .A2(new_n337_), .A3(new_n654_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G64gat), .B1(new_n740_), .B2(new_n562_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT48), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n738_), .A2(new_n747_), .A3(new_n658_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G71gat), .B1(new_n740_), .B2(new_n580_), .ZN(new_n749_));
  XOR2_X1   g548(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n738_), .A2(new_n753_), .A3(new_n533_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G78gat), .B1(new_n740_), .B2(new_n692_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1335gat));
  AND2_X1   g556(.A1(new_n737_), .A2(new_n672_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n552_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n613_), .A2(new_n634_), .A3(new_n363_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n686_), .A2(new_n697_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n763_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n551_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT108), .Z(new_n768_));
  AOI21_X1  g567(.A(new_n759_), .B1(new_n766_), .B2(new_n768_), .ZN(G1336gat));
  NAND3_X1  g568(.A1(new_n758_), .A2(new_n208_), .A3(new_n654_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n766_), .A2(new_n654_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n208_), .ZN(G1337gat));
  AOI21_X1  g571(.A(new_n240_), .B1(new_n766_), .B2(new_n658_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n418_), .A2(new_n220_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n758_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT51), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n580_), .B(new_n761_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n778_), .B(new_n775_), .C1(new_n779_), .C2(new_n240_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1338gat));
  NOR2_X1   g580(.A1(new_n692_), .A2(G106gat), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n735_), .A2(new_n736_), .A3(new_n672_), .A4(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT109), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n761_), .A2(new_n692_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n221_), .B1(new_n762_), .B2(new_n785_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n786_), .A2(KEYINPUT52), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(KEYINPUT52), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1339gat));
  NAND2_X1  g590(.A1(new_n687_), .A2(new_n552_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(KEYINPUT59), .ZN(new_n793_));
  NOR4_X1   g592(.A1(new_n309_), .A2(new_n634_), .A3(new_n612_), .A4(new_n364_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT54), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n595_), .A2(new_n600_), .A3(new_n606_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n633_), .A2(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n267_), .A2(new_n269_), .A3(new_n584_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n593_), .B1(new_n599_), .B2(KEYINPUT12), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n596_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT12), .B1(new_n247_), .B2(new_n350_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n597_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n805_), .A2(KEYINPUT55), .A3(new_n586_), .A4(new_n585_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n595_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT111), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n595_), .A2(new_n811_), .A3(new_n808_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n807_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT112), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n803_), .A2(new_n806_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n811_), .B1(new_n595_), .B2(new_n808_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n812_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n605_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n822_), .B(new_n606_), .C1(new_n814_), .C2(new_n819_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n800_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n615_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n616_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n629_), .B1(new_n826_), .B2(new_n614_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n827_), .A3(new_n625_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n625_), .B1(new_n618_), .B2(new_n631_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT113), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n624_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n828_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n834_), .A3(new_n608_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n797_), .B(new_n306_), .C1(new_n824_), .C2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n831_), .A2(new_n834_), .A3(new_n798_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n818_), .B1(new_n817_), .B2(new_n812_), .ZN(new_n838_));
  AND4_X1   g637(.A1(new_n818_), .A2(new_n807_), .A3(new_n812_), .A4(new_n810_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n605_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n822_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n605_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n837_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n309_), .B1(new_n843_), .B2(KEYINPUT58), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n831_), .A2(new_n834_), .A3(new_n798_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n845_), .B(KEYINPUT58), .C1(new_n821_), .C2(new_n823_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n306_), .B1(new_n824_), .B2(new_n835_), .ZN(new_n848_));
  OAI22_X1  g647(.A1(new_n844_), .A2(new_n847_), .B1(new_n848_), .B2(KEYINPUT57), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n836_), .B1(new_n849_), .B2(KEYINPUT116), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n634_), .A2(new_n798_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n835_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n671_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n797_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n855_), .B(new_n856_), .C1(new_n847_), .C2(new_n844_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n363_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n796_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI211_X1 g659(.A(KEYINPUT117), .B(new_n363_), .C1(new_n850_), .C2(new_n857_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n793_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT114), .B1(new_n844_), .B2(new_n847_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n845_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n309_), .A4(new_n846_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n848_), .A2(KEYINPUT57), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n863_), .A2(new_n868_), .A3(new_n855_), .A4(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n363_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n824_), .A2(new_n835_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n873_), .B2(new_n671_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n836_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n875_), .A2(KEYINPUT115), .A3(new_n863_), .A4(new_n868_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n795_), .B1(new_n872_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT59), .B1(new_n877_), .B2(new_n792_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n862_), .A2(new_n634_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G113gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n855_), .A2(new_n869_), .A3(new_n868_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n683_), .B1(new_n865_), .B2(new_n864_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n867_), .B1(new_n882_), .B2(new_n846_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n871_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n876_), .A3(new_n364_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n796_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n792_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OR3_X1    g687(.A1(new_n888_), .A2(G113gat), .A3(new_n633_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n880_), .A2(new_n889_), .ZN(G1340gat));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT118), .B(G120gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n613_), .B2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n886_), .A2(new_n887_), .A3(new_n894_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n862_), .A2(new_n878_), .A3(new_n612_), .A4(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n893_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n895_), .A2(KEYINPUT60), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1341gat));
  INV_X1    g698(.A(new_n888_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G127gat), .B1(new_n900_), .B2(new_n363_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n862_), .A2(new_n878_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n363_), .A2(G127gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT119), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n901_), .B1(new_n902_), .B2(new_n904_), .ZN(G1342gat));
  NAND3_X1  g704(.A1(new_n862_), .A2(new_n309_), .A3(new_n878_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(G134gat), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n888_), .A2(G134gat), .A3(new_n671_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1343gat));
  XNOR2_X1  g708(.A(KEYINPUT121), .B(G141gat), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n580_), .A2(new_n552_), .A3(new_n533_), .A4(new_n562_), .ZN(new_n912_));
  XOR2_X1   g711(.A(new_n912_), .B(KEYINPUT120), .Z(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n885_), .B2(new_n796_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n916_), .A3(new_n634_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n915_), .B2(new_n634_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n911_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n919_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n917_), .A3(new_n910_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(G1344gat));
  NAND2_X1  g722(.A1(new_n915_), .A2(new_n612_), .ZN(new_n924_));
  XOR2_X1   g723(.A(KEYINPUT123), .B(G148gat), .Z(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1345gat));
  NAND2_X1  g725(.A1(new_n915_), .A2(new_n363_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT61), .B(G155gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  NAND2_X1  g728(.A1(new_n886_), .A2(new_n913_), .ZN(new_n930_));
  OR3_X1    g729(.A1(new_n930_), .A2(G162gat), .A3(new_n671_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G162gat), .B1(new_n930_), .B2(new_n683_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n580_), .A2(new_n552_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n654_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n533_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n634_), .B(new_n936_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G169gat), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n937_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n860_), .A2(new_n861_), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n942_), .A2(new_n634_), .A3(new_n428_), .A4(new_n936_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n940_), .A2(new_n941_), .A3(new_n943_), .ZN(G1348gat));
  NAND2_X1  g743(.A1(new_n612_), .A2(G176gat), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n877_), .A2(new_n533_), .A3(new_n935_), .A4(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n942_), .A2(new_n612_), .A3(new_n936_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n429_), .ZN(G1349gat));
  NOR2_X1   g747(.A1(new_n935_), .A2(new_n364_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n886_), .A2(new_n692_), .A3(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n886_), .A2(new_n692_), .A3(new_n949_), .ZN(new_n953_));
  AOI21_X1  g752(.A(G183gat), .B1(new_n953_), .B2(KEYINPUT124), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n860_), .A2(new_n861_), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n955_), .A2(new_n533_), .A3(new_n935_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n364_), .A2(new_n381_), .ZN(new_n957_));
  AOI22_X1  g756(.A1(new_n952_), .A2(new_n954_), .B1(new_n956_), .B2(new_n957_), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n942_), .A2(new_n309_), .A3(new_n936_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(G190gat), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n942_), .A2(new_n382_), .A3(new_n306_), .A4(new_n936_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1351gat));
  NAND2_X1  g761(.A1(new_n580_), .A2(new_n689_), .ZN(new_n963_));
  XOR2_X1   g762(.A(new_n963_), .B(KEYINPUT125), .Z(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(new_n654_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n877_), .A2(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n634_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g767(.A(new_n965_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n886_), .A2(new_n969_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n970_), .A2(new_n613_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1353gat));
  AOI211_X1 g772(.A(KEYINPUT63), .B(G211gat), .C1(new_n966_), .C2(new_n363_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(KEYINPUT63), .B(G211gat), .ZN(new_n975_));
  NOR3_X1   g774(.A1(new_n970_), .A2(new_n364_), .A3(new_n975_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n974_), .A2(new_n976_), .ZN(G1354gat));
  INV_X1    g776(.A(G218gat), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n978_), .B1(new_n966_), .B2(new_n309_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n671_), .A2(G218gat), .ZN(new_n980_));
  AND3_X1   g779(.A1(new_n886_), .A2(new_n969_), .A3(new_n980_), .ZN(new_n981_));
  OAI21_X1  g780(.A(KEYINPUT127), .B1(new_n979_), .B2(new_n981_), .ZN(new_n982_));
  INV_X1    g781(.A(new_n981_), .ZN(new_n983_));
  OAI21_X1  g782(.A(G218gat), .B1(new_n970_), .B2(new_n683_), .ZN(new_n984_));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n983_), .A2(new_n984_), .A3(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n982_), .A2(new_n986_), .ZN(G1355gat));
endmodule


