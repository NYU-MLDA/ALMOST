//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n989_, new_n990_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT102), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT7), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n204_), .B(new_n208_), .C1(new_n210_), .C2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G85gat), .B(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n207_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G85gat), .ZN(new_n227_));
  INV_X1    g026(.A(G92gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT9), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT9), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(KEYINPUT9), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n226_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n233_), .A2(new_n230_), .A3(new_n229_), .A4(new_n234_), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n217_), .A2(new_n219_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G29gat), .B(G36gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G43gat), .B(G50gat), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G232gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT34), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT68), .B(KEYINPUT35), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n238_), .A2(new_n245_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n235_), .A2(new_n231_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n252_), .A2(new_n237_), .A3(new_n225_), .A4(new_n222_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n204_), .ZN(new_n254_));
  NOR3_X1   g053(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AOI211_X1 g055(.A(KEYINPUT8), .B(new_n214_), .C1(new_n256_), .C2(new_n225_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n218_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n253_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n241_), .A2(new_n244_), .A3(KEYINPUT15), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT15), .B1(new_n241_), .B2(new_n244_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n247_), .A2(new_n249_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT69), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n251_), .B(new_n263_), .C1(new_n264_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n248_), .A2(new_n250_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n245_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n264_), .B(new_n268_), .C1(new_n259_), .C2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n263_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n259_), .B2(new_n269_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n270_), .B(new_n271_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G190gat), .B(G218gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(KEYINPUT36), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n267_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT71), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n267_), .A2(new_n274_), .A3(new_n281_), .A4(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n267_), .A2(new_n274_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n277_), .B(KEYINPUT36), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT101), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT101), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n289_), .A3(new_n286_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT25), .B(G183gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G190gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT78), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT78), .B1(new_n293_), .B2(new_n294_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT23), .ZN(new_n300_));
  OR2_X1    g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT24), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(KEYINPUT24), .A3(new_n303_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n300_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT80), .B(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT22), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(G169gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT22), .B(G169gat), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n306_), .B(new_n309_), .C1(new_n310_), .C2(new_n307_), .ZN(new_n311_));
  OR2_X1    g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n300_), .A2(new_n312_), .B1(G169gat), .B2(G176gat), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n298_), .A2(new_n305_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G227gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(G15gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT30), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n314_), .A2(new_n318_), .ZN(new_n320_));
  INV_X1    g119(.A(G134gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G127gat), .ZN(new_n322_));
  INV_X1    g121(.A(G127gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G134gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G120gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G113gat), .ZN(new_n327_));
  INV_X1    g126(.A(G113gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G120gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n322_), .A2(new_n324_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT81), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT81), .B1(new_n331_), .B2(new_n332_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n319_), .A2(new_n320_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339_));
  INV_X1    g138(.A(G43gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT31), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n336_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n338_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  INV_X1    g154(.A(G141gat), .ZN(new_n356_));
  INV_X1    g155(.A(G148gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n357_), .A3(KEYINPUT3), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n353_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n351_), .A2(KEYINPUT82), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(G141gat), .A3(G148gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n362_), .A3(new_n352_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n350_), .B1(new_n359_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n356_), .A2(new_n357_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n360_), .A2(new_n362_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT1), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n333_), .A2(new_n334_), .B1(new_n364_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n359_), .A2(new_n363_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n349_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n331_), .A2(new_n332_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n370_), .A2(new_n375_), .A3(KEYINPUT4), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT94), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT94), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n370_), .A2(new_n375_), .A3(new_n378_), .A4(KEYINPUT4), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n372_), .A2(new_n373_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n335_), .A2(new_n382_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT95), .B1(new_n370_), .B2(KEYINPUT4), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n381_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n380_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n370_), .A2(new_n375_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n381_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT96), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT96), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n370_), .A2(new_n375_), .A3(new_n392_), .A4(new_n381_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT0), .B(G57gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n388_), .A2(new_n399_), .A3(new_n394_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT19), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT88), .ZN(new_n406_));
  INV_X1    g205(.A(G218gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G211gat), .ZN(new_n408_));
  INV_X1    g207(.A(G211gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G218gat), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n408_), .A2(new_n410_), .A3(KEYINPUT87), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT87), .B1(new_n408_), .B2(new_n410_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G197gat), .A2(G204gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G197gat), .A2(G204gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(KEYINPUT21), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT21), .ZN(new_n418_));
  INV_X1    g217(.A(new_n416_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n414_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n406_), .B1(new_n413_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n409_), .A2(G218gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n407_), .A2(G211gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n408_), .A2(new_n410_), .A3(KEYINPUT87), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n428_), .A2(KEYINPUT88), .A3(new_n417_), .A4(new_n420_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n422_), .A2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n419_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n426_), .A2(new_n431_), .A3(new_n427_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n426_), .A2(new_n431_), .A3(KEYINPUT89), .A4(new_n427_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n298_), .A2(new_n305_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n313_), .A2(new_n311_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT20), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n300_), .A2(new_n312_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n310_), .A2(new_n306_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n303_), .B(KEYINPUT91), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n443_), .A2(KEYINPUT92), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT92), .B1(new_n443_), .B2(new_n444_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n442_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n293_), .A2(new_n294_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n448_), .A2(new_n300_), .A3(new_n302_), .A4(new_n304_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n430_), .A2(new_n436_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n405_), .B1(new_n441_), .B2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G8gat), .B(G36gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT32), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n437_), .A2(new_n440_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n422_), .A2(new_n429_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n405_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n458_), .A2(new_n460_), .A3(KEYINPUT20), .A4(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n451_), .A2(new_n457_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT98), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT98), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n451_), .A2(new_n465_), .A3(new_n457_), .A4(new_n462_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n459_), .B2(new_n314_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n447_), .A2(new_n449_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n437_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n471_), .A3(new_n461_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT99), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n458_), .A2(new_n460_), .A3(KEYINPUT20), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n405_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT99), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n469_), .A2(new_n471_), .A3(new_n476_), .A4(new_n461_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n457_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n403_), .A2(new_n467_), .A3(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n451_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n456_), .B1(new_n451_), .B2(new_n462_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n380_), .A2(new_n387_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(KEYINPUT33), .A3(new_n399_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n402_), .A2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n390_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n380_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n389_), .A2(KEYINPUT97), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n381_), .B1(new_n389_), .B2(KEYINPUT97), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n399_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n484_), .A2(new_n486_), .A3(new_n488_), .A4(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n481_), .A2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(KEYINPUT85), .A2(G233gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(KEYINPUT85), .A2(G233gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(G228gat), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT86), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n384_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n437_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT29), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n500_), .B1(new_n459_), .B2(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n505_), .A2(new_n508_), .A3(G78gat), .ZN(new_n509_));
  AOI21_X1  g308(.A(G78gat), .B1(new_n505_), .B2(new_n508_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n207_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G78gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n507_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n501_), .B1(new_n437_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n502_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n459_), .A2(new_n515_), .A3(new_n500_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n512_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n505_), .A2(new_n508_), .A3(G78gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(G106gat), .A3(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n511_), .A2(KEYINPUT84), .A3(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT28), .B1(new_n384_), .B2(KEYINPUT29), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n372_), .A2(new_n522_), .A3(new_n506_), .A4(new_n373_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT83), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G22gat), .B(G50gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT83), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n521_), .A2(new_n527_), .A3(new_n523_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n529_), .A2(new_n530_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n533_), .A2(new_n511_), .A3(KEYINPUT84), .A4(new_n519_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n496_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n534_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n451_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT27), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n456_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n478_), .A2(new_n541_), .ZN(new_n542_));
  AND4_X1   g341(.A1(KEYINPUT20), .A2(new_n458_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n461_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n541_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n538_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT27), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n540_), .A2(new_n542_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n403_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n537_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n346_), .B1(new_n536_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n346_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n539_), .B1(new_n541_), .B2(new_n478_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT27), .B1(new_n545_), .B2(new_n538_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT100), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n540_), .A2(new_n542_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n546_), .A2(new_n547_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT100), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n552_), .B(new_n537_), .C1(new_n555_), .C2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n203_), .B(new_n292_), .C1(new_n551_), .C2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n552_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n553_), .A2(KEYINPUT100), .A3(new_n554_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n558_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n535_), .B(new_n563_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n403_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n496_), .A2(new_n535_), .B1(new_n567_), .B2(new_n548_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n568_), .B2(new_n346_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n203_), .B1(new_n569_), .B2(new_n292_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n562_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572_));
  INV_X1    g371(.A(G8gat), .ZN(new_n573_));
  NOR2_X1   g372(.A1(KEYINPUT72), .A2(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(KEYINPUT72), .A2(G1gat), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n573_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT14), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n572_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G1gat), .B(G8gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n576_), .ZN(new_n583_));
  OAI21_X1  g382(.A(G8gat), .B1(new_n583_), .B2(new_n574_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT14), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n572_), .A3(new_n580_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT73), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n587_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G57gat), .B(G64gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT11), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(KEYINPUT11), .ZN(new_n594_));
  INV_X1    g393(.A(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n591_), .A2(KEYINPUT11), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n590_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n590_), .A2(new_n599_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n600_), .A2(KEYINPUT74), .A3(new_n601_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n605_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(KEYINPUT17), .A2(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n607_), .A2(KEYINPUT17), .A3(new_n608_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT15), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n245_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n241_), .A2(new_n244_), .A3(KEYINPUT15), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT75), .B1(new_n615_), .B2(new_n587_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n586_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n580_), .B1(new_n585_), .B2(new_n572_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n262_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n245_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(new_n269_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n624_), .B1(new_n628_), .B2(new_n623_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(G113gat), .B(G141gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(G169gat), .B(G197gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT76), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT77), .B1(new_n631_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n625_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT77), .B(new_n635_), .C1(new_n638_), .C2(new_n629_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n627_), .A2(new_n630_), .A3(new_n634_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT13), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT66), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT5), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n648_), .B(new_n649_), .Z(new_n650_));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n598_), .B(new_n253_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT12), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n217_), .A2(new_n219_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n598_), .B1(new_n654_), .B2(new_n253_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT12), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n259_), .A2(new_n657_), .A3(new_n599_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n651_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n259_), .A2(new_n599_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n651_), .B1(new_n661_), .B2(new_n652_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT65), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n651_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(KEYINPUT12), .A3(new_n652_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n658_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT65), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n662_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n646_), .B(new_n650_), .C1(new_n664_), .C2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n650_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n660_), .A2(new_n671_), .A3(new_n663_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n660_), .A2(KEYINPUT65), .A3(new_n663_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n668_), .B1(new_n667_), .B2(new_n662_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n646_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n645_), .B1(new_n673_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n672_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n676_), .B2(new_n646_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n650_), .B1(new_n664_), .B2(new_n669_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT66), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n680_), .A2(KEYINPUT13), .A3(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n678_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT67), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n678_), .A2(new_n683_), .A3(KEYINPUT67), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n644_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n571_), .A2(new_n611_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n202_), .B1(new_n690_), .B2(new_n403_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n545_), .A2(new_n538_), .A3(new_n494_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT33), .B1(new_n485_), .B2(new_n399_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n401_), .A2(new_n402_), .B1(new_n479_), .B2(new_n478_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n486_), .A2(new_n694_), .B1(new_n695_), .B2(new_n467_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n550_), .B1(new_n696_), .B2(new_n537_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n346_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n537_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n697_), .A2(new_n698_), .B1(new_n699_), .B2(new_n563_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n644_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n686_), .A2(new_n687_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT37), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n287_), .B(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n611_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n701_), .A2(new_n702_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT38), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n403_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n707_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n691_), .A2(new_n711_), .A3(KEYINPUT103), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT103), .B1(new_n691_), .B2(new_n711_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1324gat));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n611_), .B(new_n644_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n564_), .A2(new_n565_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n716_), .B(new_n717_), .C1(new_n562_), .C2(new_n570_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(KEYINPUT104), .A3(G8gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT104), .B1(new_n718_), .B2(G8gat), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT39), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(G8gat), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n721_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n706_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n573_), .A3(new_n717_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n715_), .B1(new_n722_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n723_), .A2(new_n724_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n718_), .A2(KEYINPUT104), .A3(G8gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(KEYINPUT39), .A3(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n732_), .A2(KEYINPUT40), .A3(new_n725_), .A4(new_n727_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(new_n733_), .ZN(G1325gat));
  NAND3_X1  g533(.A1(new_n726_), .A2(new_n316_), .A3(new_n346_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n690_), .A2(new_n346_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT41), .B1(new_n736_), .B2(G15gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(G1326gat));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n690_), .A2(new_n537_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G22gat), .ZN(new_n742_));
  INV_X1    g541(.A(G22gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT42), .B(new_n743_), .C1(new_n690_), .C2(new_n537_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n537_), .A2(new_n743_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT105), .Z(new_n746_));
  OAI22_X1  g545(.A1(new_n742_), .A2(new_n744_), .B1(new_n706_), .B2(new_n746_), .ZN(G1327gat));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n748_));
  INV_X1    g547(.A(new_n704_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n700_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n569_), .A2(KEYINPUT43), .A3(new_n704_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n750_), .A2(new_n611_), .A3(new_n688_), .A4(new_n751_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n611_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n569_), .A2(new_n704_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n748_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n757_), .A2(KEYINPUT44), .A3(new_n688_), .A4(new_n751_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n754_), .A2(new_n758_), .A3(G29gat), .A4(new_n403_), .ZN(new_n759_));
  INV_X1    g558(.A(G29gat), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n292_), .A2(new_n755_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n701_), .A2(new_n702_), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n762_), .B2(new_n549_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n759_), .A2(new_n763_), .ZN(G1328gat));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n717_), .A3(new_n758_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G36gat), .ZN(new_n766_));
  INV_X1    g565(.A(new_n717_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n767_), .A2(G36gat), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n762_), .A2(KEYINPUT45), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT45), .B1(new_n762_), .B2(new_n768_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n766_), .A2(new_n771_), .A3(KEYINPUT46), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1329gat));
  NAND4_X1  g575(.A1(new_n754_), .A2(new_n758_), .A3(G43gat), .A4(new_n346_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n340_), .B1(new_n762_), .B2(new_n698_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(G1330gat));
  NAND4_X1  g580(.A1(new_n754_), .A2(new_n758_), .A3(G50gat), .A4(new_n537_), .ZN(new_n782_));
  INV_X1    g581(.A(G50gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n762_), .B2(new_n535_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1331gat));
  NOR3_X1   g584(.A1(new_n700_), .A2(new_n702_), .A3(new_n643_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(new_n705_), .ZN(new_n787_));
  INV_X1    g586(.A(G57gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n403_), .ZN(new_n789_));
  NOR4_X1   g588(.A1(new_n571_), .A2(new_n611_), .A3(new_n702_), .A4(new_n643_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n790_), .A2(new_n403_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n791_), .B2(new_n788_), .ZN(G1332gat));
  INV_X1    g591(.A(G64gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n793_), .A3(new_n717_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT48), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n790_), .A2(new_n717_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(G64gat), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT48), .B(new_n793_), .C1(new_n790_), .C2(new_n717_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(G1333gat));
  NOR2_X1   g598(.A1(new_n698_), .A2(G71gat), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT109), .Z(new_n801_));
  NAND2_X1  g600(.A1(new_n787_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n790_), .A2(new_n346_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n804_));
  AND3_X1   g603(.A1(new_n803_), .A2(G71gat), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(G71gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(G1334gat));
  NAND3_X1  g606(.A1(new_n787_), .A2(new_n512_), .A3(new_n537_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n790_), .A2(new_n537_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(G78gat), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT50), .B(new_n512_), .C1(new_n790_), .C2(new_n537_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(G1335gat));
  AND2_X1   g612(.A1(new_n786_), .A2(new_n761_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n227_), .A3(new_n403_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n702_), .A2(new_n643_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n757_), .A2(new_n751_), .A3(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n817_), .A2(new_n403_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n815_), .B1(new_n818_), .B2(new_n227_), .ZN(G1336gat));
  NAND2_X1  g618(.A1(new_n786_), .A2(new_n761_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n228_), .B1(new_n820_), .B2(new_n767_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n821_), .A2(KEYINPUT110), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(KEYINPUT110), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n767_), .A2(new_n228_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n822_), .A2(new_n823_), .B1(new_n817_), .B2(new_n824_), .ZN(G1337gat));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n346_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n814_), .A2(new_n826_), .A3(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT112), .B1(new_n820_), .B2(new_n827_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n757_), .A2(new_n346_), .A3(new_n751_), .A4(new_n816_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n832_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT111), .B1(new_n832_), .B2(G99gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n831_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT51), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n831_), .B(new_n837_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1338gat));
  NAND3_X1  g638(.A1(new_n814_), .A2(new_n207_), .A3(new_n537_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n757_), .A2(new_n537_), .A3(new_n751_), .A4(new_n816_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(new_n842_), .A3(G106gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n841_), .B2(G106gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n840_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT53), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n840_), .B(new_n847_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1339gat));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n622_), .A2(G229gat), .A3(G233gat), .A4(new_n623_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n628_), .A2(new_n623_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n634_), .B1(new_n852_), .B2(new_n624_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n672_), .A2(new_n640_), .A3(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n667_), .B(KEYINPUT55), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n666_), .A2(new_n658_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n651_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n650_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n859_), .B2(KEYINPUT56), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n660_), .A2(KEYINPUT55), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n667_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n858_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n861_), .B1(new_n866_), .B2(new_n650_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n850_), .B1(new_n860_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n859_), .A2(KEYINPUT56), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n861_), .A3(new_n650_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(KEYINPUT58), .A4(new_n855_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n868_), .A2(new_n704_), .A3(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n640_), .B(new_n854_), .C1(new_n673_), .C2(new_n677_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n672_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI22_X1  g675(.A1(new_n865_), .A2(new_n671_), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT114), .B(new_n672_), .C1(new_n636_), .C2(new_n641_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n650_), .B(new_n879_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .A4(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n291_), .B1(new_n873_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n872_), .B1(new_n882_), .B2(KEYINPUT57), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n884_), .B(new_n291_), .C1(new_n873_), .C2(new_n881_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n611_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n611_), .A2(new_n643_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n678_), .A2(new_n683_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT113), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n678_), .A2(new_n683_), .A3(new_n888_), .A4(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n887_), .B1(new_n893_), .B2(new_n749_), .ZN(new_n894_));
  AOI211_X1 g693(.A(KEYINPUT54), .B(new_n704_), .C1(new_n890_), .C2(new_n892_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n886_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n699_), .A2(new_n403_), .A3(new_n346_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n643_), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n328_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT116), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n901_), .A3(new_n328_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n896_), .A2(KEYINPUT59), .A3(new_n897_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT59), .B1(new_n896_), .B2(new_n897_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n904_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n896_), .A2(new_n897_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(KEYINPUT117), .A3(new_n905_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n644_), .A2(new_n328_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n903_), .B1(new_n913_), .B2(new_n914_), .ZN(G1340gat));
  INV_X1    g714(.A(new_n909_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n326_), .B1(new_n702_), .B2(KEYINPUT60), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n916_), .B(new_n917_), .C1(KEYINPUT60), .C2(new_n326_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n702_), .B1(new_n911_), .B2(new_n905_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n326_), .ZN(G1341gat));
  AOI21_X1  g719(.A(G127gat), .B1(new_n916_), .B2(new_n755_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n611_), .A2(new_n323_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n913_), .B2(new_n922_), .ZN(G1342gat));
  AOI21_X1  g722(.A(G134gat), .B1(new_n916_), .B2(new_n291_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n704_), .A2(G134gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT118), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n913_), .B2(new_n926_), .ZN(G1343gat));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n767_), .A2(new_n403_), .A3(new_n537_), .A4(new_n698_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT119), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n896_), .A2(new_n928_), .A3(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n928_), .B1(new_n896_), .B2(new_n930_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n643_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g733(.A(new_n702_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g736(.A(new_n755_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT61), .B(G155gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1346gat));
  OAI21_X1  g739(.A(new_n704_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(G162gat), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n292_), .A2(G162gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n942_), .A2(new_n944_), .ZN(G1347gat));
  NOR3_X1   g744(.A1(new_n767_), .A2(new_n537_), .A3(new_n552_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n896_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n643_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(G169gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n951_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n949_), .A2(G169gat), .A3(new_n953_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n948_), .A2(new_n310_), .A3(new_n643_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n952_), .A2(new_n954_), .A3(new_n955_), .ZN(G1348gat));
  NAND2_X1  g755(.A1(new_n948_), .A2(new_n935_), .ZN(new_n957_));
  INV_X1    g756(.A(G176gat), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n959_), .B1(new_n306_), .B2(new_n957_), .ZN(G1349gat));
  INV_X1    g759(.A(G183gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(new_n947_), .B2(new_n611_), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n963_));
  INV_X1    g762(.A(new_n293_), .ZN(new_n964_));
  NAND4_X1  g763(.A1(new_n896_), .A2(new_n964_), .A3(new_n755_), .A4(new_n946_), .ZN(new_n965_));
  AND3_X1   g764(.A1(new_n962_), .A2(new_n963_), .A3(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n963_), .B1(new_n962_), .B2(new_n965_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n966_), .A2(new_n967_), .ZN(G1350gat));
  OAI21_X1  g767(.A(G190gat), .B1(new_n947_), .B2(new_n749_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n291_), .A2(new_n294_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n969_), .B1(new_n947_), .B2(new_n970_), .ZN(G1351gat));
  AOI21_X1  g770(.A(KEYINPUT123), .B1(new_n567_), .B2(new_n698_), .ZN(new_n972_));
  AND3_X1   g771(.A1(new_n567_), .A2(KEYINPUT123), .A3(new_n698_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n767_), .A2(new_n972_), .A3(new_n973_), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n896_), .A2(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(new_n643_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n935_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g778(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n980_), .A2(KEYINPUT125), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n611_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n982_));
  XNOR2_X1  g781(.A(new_n982_), .B(KEYINPUT124), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n981_), .B1(new_n975_), .B2(new_n983_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n980_), .A2(KEYINPUT125), .ZN(new_n985_));
  XOR2_X1   g784(.A(new_n985_), .B(KEYINPUT126), .Z(new_n986_));
  XNOR2_X1  g785(.A(new_n984_), .B(new_n986_), .ZN(G1354gat));
  INV_X1    g786(.A(new_n975_), .ZN(new_n988_));
  OAI21_X1  g787(.A(G218gat), .B1(new_n988_), .B2(new_n749_), .ZN(new_n989_));
  NAND3_X1  g788(.A1(new_n975_), .A2(new_n407_), .A3(new_n291_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n989_), .A2(new_n990_), .ZN(G1355gat));
endmodule


