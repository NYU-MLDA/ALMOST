//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G85gat), .B(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT9), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G85gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(G92gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n209_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT65), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AOI211_X1 g023(.A(new_n207_), .B(new_n220_), .C1(new_n224_), .C2(new_n214_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n204_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n212_), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n221_), .B(new_n229_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n207_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n226_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT67), .B1(new_n225_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n220_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n211_), .A2(new_n213_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(new_n221_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n233_), .B(new_n236_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n207_), .B1(new_n224_), .B2(new_n214_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n239_), .B(new_n240_), .C1(new_n241_), .C2(new_n226_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n218_), .B1(new_n235_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G78gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(KEYINPUT11), .B2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n244_), .A3(KEYINPUT11), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT12), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n233_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n226_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n218_), .B1(new_n255_), .B2(new_n239_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(new_n250_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n256_), .B2(new_n250_), .ZN(new_n259_));
  OAI221_X1 g058(.A(new_n202_), .B1(new_n243_), .B2(new_n252_), .C1(new_n257_), .C2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n202_), .B1(new_n257_), .B2(KEYINPUT66), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n239_), .B1(new_n241_), .B2(new_n226_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n209_), .A2(new_n217_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n251_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n250_), .A3(new_n263_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G120gat), .B(G148gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT5), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G176gat), .B(G204gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n260_), .A2(new_n269_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT68), .ZN(new_n276_));
  INV_X1    g075(.A(new_n242_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n240_), .B1(new_n255_), .B2(new_n239_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n263_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n252_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n267_), .A2(KEYINPUT12), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n279_), .A2(new_n280_), .B1(new_n281_), .B2(new_n265_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n282_), .A2(new_n202_), .B1(new_n268_), .B2(new_n261_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n274_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n276_), .A2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n283_), .A2(new_n274_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT13), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(KEYINPUT13), .A3(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT15), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G15gat), .B(G22gat), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n293_), .B(new_n294_), .Z(new_n305_));
  OR2_X1    g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT77), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n303_), .B(new_n305_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(G229gat), .A3(G233gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT79), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G113gat), .B(G141gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT78), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G169gat), .B(G197gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT79), .B1(new_n309_), .B2(new_n311_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n292_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G71gat), .B(G99gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G43gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT84), .B(G15gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT80), .B(G183gat), .ZN(new_n332_));
  INV_X1    g131(.A(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G183gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT23), .B1(new_n335_), .B2(new_n333_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT82), .B(G169gat), .ZN(new_n342_));
  OR2_X1    g141(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n343_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n340_), .A2(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n334_), .A2(new_n339_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT83), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT81), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n338_), .A2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n338_), .A2(new_n349_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n336_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G169gat), .ZN(new_n353_));
  INV_X1    g152(.A(G176gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(KEYINPUT24), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(KEYINPUT24), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n335_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n332_), .B2(new_n360_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G190gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n359_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n346_), .A2(new_n348_), .B1(new_n352_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT30), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n331_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n367_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G113gat), .B(G120gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(KEYINPUT86), .ZN(new_n374_));
  INV_X1    g173(.A(G134gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G127gat), .ZN(new_n376_));
  INV_X1    g175(.A(G127gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G134gat), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n376_), .A2(new_n378_), .A3(KEYINPUT86), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n372_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n378_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n373_), .A2(KEYINPUT86), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(new_n371_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n386_), .B(KEYINPUT31), .Z(new_n387_));
  OR2_X1    g186(.A1(new_n370_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n370_), .A2(new_n387_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT87), .B1(new_n391_), .B2(KEYINPUT1), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT1), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(G155gat), .A4(G162gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(KEYINPUT1), .ZN(new_n396_));
  OR2_X1    g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n392_), .A2(new_n395_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G141gat), .B(G148gat), .Z(new_n399_));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400_));
  INV_X1    g199(.A(G141gat), .ZN(new_n401_));
  INV_X1    g200(.A(G148gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n403_), .A2(new_n406_), .A3(new_n407_), .A4(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n397_), .A2(new_n391_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n398_), .A2(new_n399_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(KEYINPUT28), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(KEYINPUT28), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G22gat), .B(G50gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(G197gat), .A2(G204gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G197gat), .A2(G204gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(KEYINPUT21), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G211gat), .B(G218gat), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428_));
  XOR2_X1   g227(.A(G197gat), .B(G204gat), .Z(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n429_), .B2(KEYINPUT21), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n422_), .A2(new_n423_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT21), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT90), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n424_), .A2(KEYINPUT89), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n422_), .A2(new_n436_), .A3(KEYINPUT21), .A4(new_n423_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n426_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n434_), .A2(new_n438_), .A3(KEYINPUT91), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT91), .B1(new_n434_), .B2(new_n438_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n427_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442_));
  INV_X1    g241(.A(G228gat), .ZN(new_n443_));
  INV_X1    g242(.A(G233gat), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT92), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n442_), .B(new_n445_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n398_), .A2(new_n399_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n409_), .A2(new_n410_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT29), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n446_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n441_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n442_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n441_), .A2(new_n456_), .B1(G228gat), .B2(G233gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(G78gat), .B(G106gat), .Z(new_n458_));
  NOR3_X1   g257(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n458_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n434_), .A2(new_n438_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n434_), .A2(new_n438_), .A3(KEYINPUT91), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n463_), .A2(new_n464_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n465_));
  OAI22_X1  g264(.A1(new_n465_), .A2(new_n455_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n460_), .B1(new_n466_), .B2(new_n453_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n421_), .B1(new_n459_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n458_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n453_), .A3(new_n460_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n420_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n386_), .A2(new_n449_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n411_), .A2(new_n385_), .A3(new_n380_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(KEYINPUT4), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G225gat), .A2(G233gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n474_), .B(new_n476_), .C1(KEYINPUT4), .C2(new_n472_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G29gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G85gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT0), .B(G57gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n474_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n476_), .B1(new_n472_), .B2(KEYINPUT4), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n483_), .B(new_n478_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n468_), .A2(new_n471_), .A3(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n346_), .A2(new_n348_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n364_), .A2(new_n352_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n441_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G226gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT25), .B(G183gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n363_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n339_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n503_), .A2(new_n359_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n352_), .B1(G183gat), .B2(G190gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n357_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT22), .B(G169gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(new_n354_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n504_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n509_), .B(new_n427_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n510_));
  AND4_X1   g309(.A1(KEYINPUT20), .A2(new_n496_), .A3(new_n500_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT20), .ZN(new_n512_));
  INV_X1    g311(.A(new_n509_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n441_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n465_), .A2(new_n365_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n500_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G8gat), .B(G36gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT18), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G64gat), .B(G92gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n511_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n514_), .A2(new_n515_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n499_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n512_), .B1(new_n465_), .B2(new_n509_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n500_), .A3(new_n496_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n520_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n492_), .B1(new_n522_), .B2(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n514_), .A2(new_n500_), .A3(new_n515_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n500_), .B1(new_n525_), .B2(new_n496_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n521_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n526_), .A3(new_n520_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT27), .A3(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n490_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n520_), .A2(KEYINPUT32), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n524_), .A2(new_n526_), .A3(new_n535_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n485_), .A2(new_n488_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n521_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n472_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n484_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n472_), .A2(KEYINPUT4), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(new_n476_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n545_), .B2(new_n474_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n488_), .A2(KEYINPUT33), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT33), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n477_), .A2(new_n548_), .A3(new_n483_), .A4(new_n478_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n546_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n532_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n540_), .A2(new_n551_), .B1(new_n471_), .B2(new_n468_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n534_), .B1(new_n552_), .B2(KEYINPUT94), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n540_), .A2(new_n551_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n468_), .A2(new_n471_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n554_), .A2(KEYINPUT94), .A3(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n390_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n539_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n528_), .A2(new_n533_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n555_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n325_), .B1(new_n557_), .B2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G190gat), .B(G218gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT71), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT70), .B1(new_n264_), .B2(new_n305_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT70), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n256_), .A2(new_n576_), .A3(new_n295_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n572_), .A2(new_n573_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n279_), .A2(new_n296_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n569_), .B(new_n570_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n569_), .B(KEYINPUT72), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n590_), .A3(KEYINPUT37), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT37), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n583_), .B(new_n587_), .C1(new_n589_), .C2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n303_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n250_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT17), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n597_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT75), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n602_), .A2(new_n603_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n597_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n594_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT76), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n563_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n489_), .B(KEYINPUT96), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n298_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n588_), .B(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n557_), .B2(new_n562_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n325_), .A2(new_n611_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n298_), .B1(new_n624_), .B2(new_n539_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n619_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n626_), .B1(new_n618_), .B2(new_n617_), .ZN(G1324gat));
  NAND3_X1  g426(.A1(new_n615_), .A2(new_n299_), .A3(new_n559_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n622_), .A2(new_n559_), .A3(new_n623_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n630_), .A3(G8gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n629_), .B2(G8gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT99), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT99), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1325gat));
  INV_X1    g438(.A(G15gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n390_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n624_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT41), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n615_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1326gat));
  INV_X1    g444(.A(G22gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n555_), .B(KEYINPUT100), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n624_), .B2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n615_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1327gat));
  NAND2_X1  g451(.A1(new_n557_), .A2(new_n562_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n621_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(new_n612_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n324_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n563_), .A2(KEYINPUT103), .A3(new_n655_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(G29gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n539_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n325_), .A2(new_n612_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  INV_X1    g463(.A(new_n594_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n653_), .B2(new_n665_), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT43), .B(new_n594_), .C1(new_n557_), .C2(new_n562_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT44), .B(new_n663_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(KEYINPUT102), .A3(new_n616_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G29gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT102), .B1(new_n672_), .B2(new_n616_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n662_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n670_), .A2(new_n559_), .A3(new_n671_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(G36gat), .B1(new_n528_), .B2(new_n533_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n658_), .A2(new_n659_), .A3(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT45), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT46), .B1(new_n682_), .B2(KEYINPUT104), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  AOI211_X1 g484(.A(new_n684_), .B(new_n685_), .C1(new_n678_), .C2(new_n681_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n672_), .A2(G43gat), .A3(new_n641_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n660_), .A2(new_n641_), .ZN(new_n689_));
  INV_X1    g488(.A(G43gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n688_), .A2(KEYINPUT47), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT47), .B1(new_n688_), .B2(new_n691_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1330gat));
  AOI21_X1  g493(.A(G50gat), .B1(new_n660_), .B2(new_n647_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n560_), .A2(G50gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n672_), .B2(new_n696_), .ZN(G1331gat));
  AND4_X1   g496(.A1(new_n323_), .A2(new_n622_), .A3(new_n292_), .A4(new_n612_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(G57gat), .A3(new_n539_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT106), .ZN(new_n700_));
  INV_X1    g499(.A(G57gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n292_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n653_), .A2(new_n323_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n653_), .A2(KEYINPUT105), .A3(new_n323_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n700_), .B1(new_n701_), .B2(new_n708_), .ZN(G1332gat));
  INV_X1    g508(.A(G64gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n698_), .B2(new_n559_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT48), .Z(new_n712_));
  NAND2_X1  g511(.A1(new_n707_), .A2(new_n614_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n559_), .A2(new_n710_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(G1333gat));
  NAND2_X1  g514(.A1(new_n698_), .A2(new_n641_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G71gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT107), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT49), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n717_), .B(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT49), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n713_), .A2(G71gat), .A3(new_n390_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n723_), .A3(new_n724_), .ZN(G1334gat));
  INV_X1    g524(.A(G78gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n698_), .B2(new_n647_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND2_X1  g527(.A1(new_n647_), .A2(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n713_), .B2(new_n729_), .ZN(G1335gat));
  NAND3_X1  g529(.A1(new_n292_), .A2(new_n323_), .A3(new_n611_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT109), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n733_), .A2(new_n489_), .A3(new_n215_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n705_), .A2(new_n616_), .A3(new_n655_), .A4(new_n706_), .ZN(new_n735_));
  INV_X1    g534(.A(G85gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT108), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT108), .B1(new_n735_), .B2(new_n736_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n734_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(G1336gat));
  AOI21_X1  g541(.A(new_n733_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n743_));
  INV_X1    g542(.A(G92gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n705_), .A2(new_n655_), .A3(new_n706_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n559_), .A2(new_n744_), .ZN(new_n746_));
  OAI22_X1  g545(.A1(new_n743_), .A2(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(G1337gat));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n641_), .A2(new_n203_), .A3(new_n205_), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n745_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n745_), .B2(new_n749_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G99gat), .B1(new_n733_), .B2(new_n390_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1338gat));
  XNOR2_X1  g556(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n555_), .A2(G106gat), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n745_), .A2(KEYINPUT113), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT113), .B1(new_n745_), .B2(new_n761_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n732_), .B(new_n560_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G106gat), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n759_), .B1(new_n764_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n762_), .A2(new_n763_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n758_), .C1(new_n768_), .C2(new_n767_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n611_), .B1(new_n593_), .B2(new_n591_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n702_), .A2(new_n774_), .A3(new_n775_), .A4(new_n323_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n290_), .A2(new_n323_), .A3(new_n291_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT115), .B1(new_n613_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n778_), .A3(KEYINPUT54), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT115), .B(new_n780_), .C1(new_n613_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n323_), .B1(new_n276_), .B2(new_n285_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT116), .B1(new_n282_), .B2(new_n202_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI22_X1  g584(.A1(new_n259_), .A2(new_n257_), .B1(new_n243_), .B2(new_n252_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n202_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n282_), .A2(KEYINPUT55), .A3(new_n202_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n790_), .A3(new_n787_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n784_), .A2(new_n788_), .A3(new_n789_), .A4(new_n791_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n273_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n792_), .B2(new_n273_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n783_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT118), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n783_), .B(new_n798_), .C1(new_n793_), .C2(new_n795_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n308_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n304_), .A2(new_n306_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n310_), .A2(new_n308_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n318_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n319_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n804_));
  OR3_X1    g603(.A1(new_n803_), .A2(new_n804_), .A3(KEYINPUT119), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT119), .B1(new_n804_), .B2(new_n803_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n288_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n797_), .A2(new_n799_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n654_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n621_), .A2(new_n811_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n321_), .B(new_n319_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n284_), .B1(new_n283_), .B2(new_n274_), .ZN(new_n815_));
  AND4_X1   g614(.A1(new_n284_), .A2(new_n260_), .A3(new_n269_), .A4(new_n274_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n792_), .A2(new_n273_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n794_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n273_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n817_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n808_), .B1(new_n822_), .B2(new_n798_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n799_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n813_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n273_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n793_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n807_), .A2(new_n286_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT120), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n807_), .A2(new_n832_), .A3(new_n286_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n594_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n829_), .A2(new_n831_), .A3(KEYINPUT58), .A4(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n809_), .A2(KEYINPUT121), .A3(new_n813_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n812_), .A2(new_n827_), .A3(new_n838_), .A4(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n782_), .B1(new_n840_), .B2(new_n611_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n641_), .A2(new_n561_), .A3(new_n616_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n814_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n842_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n809_), .A2(KEYINPUT121), .A3(new_n813_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT121), .B1(new_n809_), .B2(new_n813_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n810_), .A2(new_n811_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n612_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT59), .B(new_n848_), .C1(new_n853_), .C2(new_n782_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT122), .B1(new_n847_), .B2(new_n854_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n323_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n845_), .B1(new_n857_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n702_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n843_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n702_), .B1(new_n847_), .B2(new_n854_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G120gat), .B1(new_n862_), .B2(new_n863_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n861_), .B1(new_n864_), .B2(new_n865_), .ZN(G1341gat));
  NAND3_X1  g665(.A1(new_n843_), .A2(new_n377_), .A3(new_n612_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n855_), .A2(new_n856_), .A3(new_n611_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n377_), .ZN(G1342gat));
  OAI211_X1 g668(.A(new_n621_), .B(new_n848_), .C1(new_n853_), .C2(new_n782_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n375_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(KEYINPUT124), .A3(new_n375_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n855_), .A2(new_n856_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n594_), .A2(new_n375_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(G1343gat));
  INV_X1    g677(.A(new_n841_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n390_), .A2(new_n560_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n616_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n880_), .A2(new_n559_), .A3(new_n881_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT125), .Z(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n323_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n401_), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n702_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n402_), .ZN(G1345gat));
  NOR2_X1   g687(.A1(new_n884_), .A2(new_n611_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT61), .B(G155gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1346gat));
  INV_X1    g690(.A(G162gat), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n884_), .A2(new_n892_), .A3(new_n594_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n884_), .B2(new_n654_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT126), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n896_), .B(new_n892_), .C1(new_n884_), .C2(new_n654_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n893_), .B1(new_n895_), .B2(new_n897_), .ZN(G1347gat));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n641_), .A2(new_n559_), .A3(new_n881_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n841_), .A2(new_n647_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n323_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n903_), .B2(new_n353_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n507_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT62), .B(G169gat), .C1(new_n902_), .C2(new_n323_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(G1348gat));
  AOI21_X1  g706(.A(G176gat), .B1(new_n901_), .B2(new_n292_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n841_), .A2(new_n560_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n900_), .A2(new_n702_), .A3(new_n354_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1349gat));
  INV_X1    g710(.A(new_n900_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n909_), .A2(new_n612_), .A3(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n611_), .A2(new_n501_), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n913_), .A2(new_n332_), .B1(new_n901_), .B2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n902_), .B2(new_n594_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n901_), .A2(new_n363_), .A3(new_n621_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1351gat));
  NAND4_X1  g717(.A1(new_n390_), .A2(new_n560_), .A3(new_n489_), .A4(new_n559_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n841_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n814_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n292_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g723(.A1(new_n841_), .A2(new_n919_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n611_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n926_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT63), .B(G211gat), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1354gat));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n920_), .B2(new_n665_), .ZN(new_n931_));
  NOR4_X1   g730(.A1(new_n841_), .A2(G218gat), .A3(new_n654_), .A4(new_n919_), .ZN(new_n932_));
  OR3_X1    g731(.A1(new_n931_), .A2(KEYINPUT127), .A3(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT127), .B1(new_n931_), .B2(new_n932_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1355gat));
endmodule


