//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  XOR2_X1   g002(.A(G8gat), .B(G36gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G64gat), .B(G92gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(G176gat), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT94), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n219_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n218_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  AOI211_X1 g028(.A(KEYINPUT94), .B(new_n227_), .C1(new_n222_), .C2(new_n225_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n217_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G218gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G211gat), .ZN(new_n233_));
  INV_X1    g032(.A(G211gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G218gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT86), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT21), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G197gat), .A2(G204gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G197gat), .A2(G204gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n238_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n233_), .A2(new_n235_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n241_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT21), .A3(new_n239_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n237_), .A2(new_n242_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n240_), .A2(new_n241_), .A3(new_n238_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n233_), .A2(new_n235_), .A3(new_n243_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n243_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT93), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n212_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n223_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n219_), .A2(new_n224_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT26), .B(G190gat), .Z(new_n262_));
  INV_X1    g061(.A(KEYINPUT92), .ZN(new_n263_));
  INV_X1    g062(.A(G183gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT25), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT25), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n266_), .A2(G183gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n263_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(G183gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(KEYINPUT25), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(KEYINPUT92), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n262_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n254_), .B1(new_n261_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(new_n260_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT24), .ZN(new_n275_));
  INV_X1    g074(.A(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n278_), .A2(new_n255_), .B1(G169gat), .B2(G176gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n271_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT92), .B1(new_n269_), .B2(new_n270_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n284_), .A3(KEYINPUT93), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n231_), .A2(new_n253_), .A3(new_n273_), .A4(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT20), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT90), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT78), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n266_), .B2(G183gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n264_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n281_), .A2(new_n269_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n256_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n295_), .A2(new_n226_), .A3(new_n278_), .A4(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n259_), .A2(new_n228_), .A3(new_n260_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n217_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  AOI211_X1 g099(.A(new_n287_), .B(new_n291_), .C1(new_n300_), .C2(new_n252_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n273_), .A2(new_n285_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n217_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n226_), .A2(new_n228_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT94), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n226_), .A2(new_n218_), .A3(new_n228_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n252_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n297_), .A2(new_n299_), .A3(new_n247_), .A4(new_n251_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT20), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT91), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT91), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n312_), .A3(KEYINPUT20), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  AOI221_X4 g113(.A(new_n208_), .B1(new_n286_), .B2(new_n301_), .C1(new_n314_), .C2(new_n291_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n291_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n301_), .A2(new_n286_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n207_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n203_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n280_), .A2(new_n284_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n252_), .A2(KEYINPUT87), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n322_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n320_), .B(new_n231_), .C1(new_n321_), .C2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n287_), .B1(new_n300_), .B2(new_n252_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n291_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n291_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n308_), .A2(new_n311_), .A3(new_n328_), .A4(new_n313_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n208_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n316_), .A2(new_n207_), .A3(new_n317_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT27), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n319_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G227gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(G15gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT30), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G71gat), .B(G99gat), .ZN(new_n340_));
  INV_X1    g139(.A(G43gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n300_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n300_), .A2(new_n342_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n339_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n345_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(new_n338_), .A3(new_n343_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT82), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G127gat), .B(G134gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G113gat), .B(G120gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n350_), .A2(new_n351_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT81), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT31), .Z(new_n356_));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n349_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n346_), .A2(new_n348_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n356_), .B1(new_n359_), .B2(KEYINPUT83), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n349_), .A2(new_n357_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(KEYINPUT1), .B2(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n364_), .A2(KEYINPUT1), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G141gat), .B(G148gat), .Z(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT2), .ZN(new_n370_));
  INV_X1    g169(.A(G141gat), .ZN(new_n371_));
  INV_X1    g170(.A(G148gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n363_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n379_), .A2(new_n364_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n369_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n354_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n369_), .B(new_n381_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(KEYINPUT4), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n388_), .A3(new_n354_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n383_), .A2(new_n386_), .A3(new_n384_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT97), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n399_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n394_), .A2(new_n402_), .A3(new_n397_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n400_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n392_), .A2(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n404_), .A2(new_n405_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(KEYINPUT99), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT99), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n392_), .A2(new_n411_), .A3(new_n406_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n416_), .B(KEYINPUT85), .Z(new_n417_));
  AND2_X1   g216(.A1(new_n252_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n382_), .A2(KEYINPUT29), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n321_), .A2(new_n323_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n421_), .A2(new_n419_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n415_), .B(new_n420_), .C1(new_n422_), .C2(new_n417_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n415_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n417_), .B1(new_n421_), .B2(new_n419_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n420_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT28), .B1(new_n382_), .B2(KEYINPUT29), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n367_), .A2(new_n368_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G22gat), .B(G50gat), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n428_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n434_), .A2(new_n435_), .A3(KEYINPUT84), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n423_), .B(new_n427_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n424_), .A2(KEYINPUT88), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n420_), .B(new_n442_), .C1(new_n422_), .C2(new_n417_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n436_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n440_), .A2(new_n445_), .ZN(new_n446_));
  NOR4_X1   g245(.A1(new_n334_), .A2(new_n362_), .A3(new_n414_), .A4(new_n446_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n440_), .A2(new_n445_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n319_), .A3(new_n333_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n207_), .A2(KEYINPUT32), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n330_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n316_), .A2(new_n450_), .A3(new_n317_), .ZN(new_n453_));
  AND4_X1   g252(.A1(new_n412_), .A2(new_n452_), .A3(new_n410_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n409_), .A2(KEYINPUT33), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n408_), .A2(new_n390_), .A3(new_n456_), .A4(new_n391_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n385_), .A2(new_n386_), .A3(new_n389_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n383_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n406_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT98), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n459_), .A2(KEYINPUT98), .A3(new_n406_), .A4(new_n460_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n231_), .A2(new_n273_), .A3(new_n285_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n252_), .A2(new_n467_), .B1(new_n310_), .B2(KEYINPUT91), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n328_), .B1(new_n468_), .B2(new_n313_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n317_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n208_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n332_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT95), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n466_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(KEYINPUT95), .A3(new_n332_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n454_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n449_), .B1(new_n476_), .B2(new_n446_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n447_), .B1(new_n477_), .B2(new_n362_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G15gat), .B(G22gat), .ZN(new_n479_));
  INV_X1    g278(.A(G8gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G8gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G71gat), .B(G78gat), .Z(new_n486_));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n486_), .B(new_n487_), .C1(KEYINPUT11), .C2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G64gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G57gat), .ZN(new_n491_));
  INV_X1    g290(.A(G57gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G64gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT11), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G71gat), .B(G78gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT67), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n489_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n489_), .B2(new_n496_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G231gat), .A2(G233gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(new_n501_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT70), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n500_), .A2(new_n501_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(new_n502_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n485_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT70), .B1(new_n503_), .B2(new_n504_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n506_), .A3(new_n502_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n484_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT72), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT72), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n509_), .A2(new_n510_), .A3(new_n516_), .A4(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G127gat), .B(G155gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT16), .ZN(new_n520_));
  XOR2_X1   g319(.A(G183gat), .B(G211gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT17), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n509_), .A2(new_n524_), .A3(new_n513_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n525_), .B2(new_n522_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n518_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n518_), .A2(new_n526_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G85gat), .A2(G92gat), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT7), .ZN(new_n537_));
  INV_X1    g336(.A(G99gat), .ZN(new_n538_));
  INV_X1    g337(.A(G106gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n533_), .B1(new_n536_), .B2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT8), .B1(new_n533_), .B2(KEYINPUT66), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OAI221_X1 g344(.A(new_n533_), .B1(KEYINPUT66), .B2(KEYINPUT8), .C1(new_n536_), .C2(new_n542_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n531_), .A2(KEYINPUT9), .A3(new_n532_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT64), .B(G85gat), .ZN(new_n549_));
  INV_X1    g348(.A(G92gat), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT9), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n548_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT65), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n548_), .B(new_n554_), .C1(new_n549_), .C2(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT10), .B(G99gat), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n539_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n534_), .B(KEYINPUT6), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n547_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G29gat), .B(G36gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT15), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n547_), .A2(new_n566_), .A3(new_n562_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT34), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT35), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n572_), .A2(new_n573_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(new_n576_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n577_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n580_), .B(KEYINPUT36), .Z(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n577_), .B2(new_n582_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT103), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n563_), .A2(new_n500_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT68), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n545_), .A2(new_n546_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n560_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n594_));
  OAI22_X1  g393(.A1(new_n593_), .A2(new_n594_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n596_), .B(new_n598_), .C1(new_n592_), .C2(new_n591_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT69), .B1(new_n595_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n563_), .A2(new_n500_), .A3(new_n602_), .A4(KEYINPUT12), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT12), .B1(new_n563_), .B2(new_n500_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n595_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n606_), .A3(new_n597_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n599_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT5), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n610_), .B(new_n611_), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n612_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n599_), .A2(new_n607_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n590_), .B1(new_n614_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT77), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT74), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n566_), .B(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n484_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n566_), .B(KEYINPUT74), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n485_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n621_), .B2(new_n484_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n567_), .A2(new_n485_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT76), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G169gat), .B(G197gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n619_), .B1(new_n632_), .B2(new_n637_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n625_), .A2(new_n627_), .B1(new_n630_), .B2(new_n629_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(KEYINPUT77), .A3(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT75), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n632_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(KEYINPUT75), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n637_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n613_), .A2(KEYINPUT13), .A3(new_n616_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n618_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  NOR4_X1   g447(.A1(new_n478_), .A2(new_n530_), .A3(new_n589_), .A4(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n202_), .B1(new_n649_), .B2(new_n414_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n583_), .A2(new_n586_), .A3(KEYINPUT37), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT37), .B1(new_n583_), .B2(new_n586_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT73), .Z(new_n655_));
  NAND2_X1  g454(.A1(new_n618_), .A2(new_n647_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n646_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n478_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT100), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n659_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n413_), .B(KEYINPUT101), .Z(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(G1gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n661_), .A2(new_n664_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n650_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n661_), .A2(KEYINPUT38), .A3(new_n664_), .A4(new_n667_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(KEYINPUT102), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(KEYINPUT102), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(G1324gat));
  AOI21_X1  g473(.A(new_n480_), .B1(new_n649_), .B2(new_n334_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT39), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n661_), .A2(new_n664_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n334_), .A2(new_n480_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n676_), .B(KEYINPUT40), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1325gat));
  INV_X1    g482(.A(new_n362_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n660_), .A2(new_n336_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n336_), .B1(new_n649_), .B2(new_n684_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT41), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n649_), .A2(new_n446_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G22gat), .ZN(new_n690_));
  XOR2_X1   g489(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n446_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(G22gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n662_), .B2(new_n694_), .ZN(G1327gat));
  NAND2_X1  g494(.A1(new_n530_), .A2(new_n589_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n656_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(new_n659_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n414_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n529_), .A2(new_n648_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n703_));
  NAND2_X1  g502(.A1(new_n651_), .A2(new_n652_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n478_), .B2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n473_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n458_), .A2(new_n465_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n475_), .A3(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n414_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n446_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n449_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n362_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n447_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n653_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n702_), .B1(new_n705_), .B2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n700_), .B1(new_n717_), .B2(KEYINPUT44), .ZN(new_n718_));
  INV_X1    g517(.A(new_n703_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n714_), .B2(new_n653_), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT43), .B(new_n704_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n701_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(KEYINPUT106), .A3(new_n723_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n718_), .A2(new_n724_), .B1(KEYINPUT44), .B2(new_n717_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n665_), .A2(G29gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n699_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  XNOR2_X1  g526(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT44), .B(new_n701_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n334_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n718_), .B2(new_n724_), .ZN(new_n732_));
  INV_X1    g531(.A(G36gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n730_), .A2(new_n334_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n717_), .A2(new_n700_), .A3(KEYINPUT44), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n722_), .B2(new_n723_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n734_), .A2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n697_), .A2(new_n733_), .A3(new_n334_), .A4(new_n659_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n728_), .B1(new_n740_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n728_), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n743_), .B(new_n746_), .C1(new_n734_), .C2(new_n739_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1329gat));
  AOI21_X1  g547(.A(G43gat), .B1(new_n698_), .B2(new_n684_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n362_), .A2(new_n341_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n725_), .B2(new_n750_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT47), .Z(G1330gat));
  NAND2_X1  g551(.A1(new_n725_), .A2(new_n446_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n693_), .A2(G50gat), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n753_), .A2(G50gat), .B1(new_n698_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(G1331gat));
  INV_X1    g556(.A(new_n656_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n655_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n478_), .A2(new_n646_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT111), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n763_), .A3(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G57gat), .B1(new_n766_), .B2(new_n665_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n758_), .A2(new_n646_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n768_), .A2(new_n714_), .A3(new_n529_), .A4(new_n588_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT112), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(G57gat), .A3(new_n414_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n771_), .A2(new_n772_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n767_), .A2(new_n773_), .A3(new_n774_), .ZN(G1332gat));
  NAND3_X1  g574(.A1(new_n766_), .A2(new_n490_), .A3(new_n334_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n490_), .B1(new_n770_), .B2(new_n334_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT48), .Z(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n766_), .A2(new_n780_), .A3(new_n684_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n770_), .B2(new_n684_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT49), .Z(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1334gat));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n770_), .A2(new_n446_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(G78gat), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n785_), .A3(G78gat), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n693_), .A2(G78gat), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI22_X1  g589(.A1(new_n787_), .A2(new_n788_), .B1(new_n765_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI221_X1 g592(.A(KEYINPUT114), .B1(new_n765_), .B2(new_n790_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1335gat));
  NOR4_X1   g594(.A1(new_n696_), .A2(new_n478_), .A3(new_n646_), .A4(new_n758_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G85gat), .B1(new_n796_), .B2(new_n665_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n529_), .A2(new_n758_), .A3(new_n646_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n798_), .A2(KEYINPUT115), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(KEYINPUT115), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n799_), .A2(new_n800_), .B1(new_n705_), .B2(new_n716_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n413_), .A2(new_n549_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT116), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n797_), .B1(new_n801_), .B2(new_n803_), .ZN(G1336gat));
  NAND3_X1  g603(.A1(new_n796_), .A2(new_n550_), .A3(new_n334_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n801_), .A2(new_n334_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n550_), .ZN(G1337gat));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n796_), .A2(new_n684_), .A3(new_n557_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n801_), .A2(new_n684_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n808_), .B(new_n809_), .C1(new_n810_), .C2(G99gat), .ZN(new_n811_));
  XOR2_X1   g610(.A(new_n811_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g611(.A1(new_n796_), .A2(new_n539_), .A3(new_n446_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n801_), .A2(new_n446_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(G106gat), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT52), .B(new_n539_), .C1(new_n801_), .C2(new_n446_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n618_), .A2(new_n658_), .A3(new_n647_), .ZN(new_n821_));
  AND4_X1   g620(.A1(new_n820_), .A2(new_n529_), .A3(new_n821_), .A4(new_n704_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n820_), .B1(new_n654_), .B2(new_n821_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n646_), .A2(new_n616_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n597_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n607_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n604_), .A2(new_n606_), .A3(KEYINPUT55), .A4(new_n597_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n612_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n612_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n825_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n625_), .A2(new_n626_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n637_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n627_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT118), .B1(new_n839_), .B2(new_n636_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n622_), .A2(new_n630_), .A3(new_n627_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n639_), .A2(KEYINPUT77), .A3(new_n636_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT77), .B1(new_n639_), .B2(new_n636_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n641_), .A2(KEYINPUT119), .A3(new_n842_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n847_), .A2(new_n848_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT57), .B(new_n588_), .C1(new_n835_), .C2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n588_), .B1(new_n835_), .B2(new_n849_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n849_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT56), .B1(new_n830_), .B2(new_n612_), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n832_), .B(new_n615_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n859_), .B2(new_n825_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n588_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n847_), .A2(new_n848_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n616_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n859_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n833_), .A2(new_n834_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n866_), .A2(KEYINPUT58), .A3(new_n616_), .A4(new_n863_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n867_), .A3(new_n653_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n852_), .A2(new_n855_), .A3(new_n861_), .A4(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n824_), .B1(new_n869_), .B2(new_n530_), .ZN(new_n870_));
  OR4_X1    g669(.A1(new_n446_), .A2(new_n666_), .A3(new_n334_), .A4(new_n362_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT121), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G113gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n646_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n869_), .A2(new_n530_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n824_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT59), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n872_), .A3(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n870_), .B2(new_n873_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n882_), .A2(new_n885_), .A3(new_n646_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n876_), .B1(new_n886_), .B2(new_n875_), .ZN(G1340gat));
  INV_X1    g686(.A(G120gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n758_), .B2(KEYINPUT60), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n874_), .B(new_n889_), .C1(KEYINPUT60), .C2(new_n888_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n882_), .A2(new_n885_), .A3(new_n656_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n888_), .ZN(G1341gat));
  NAND3_X1  g691(.A1(new_n882_), .A2(new_n885_), .A3(new_n529_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G127gat), .ZN(new_n894_));
  INV_X1    g693(.A(G127gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n874_), .A2(new_n895_), .A3(new_n529_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT123), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n894_), .A2(new_n899_), .A3(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1342gat));
  NOR3_X1   g700(.A1(new_n870_), .A2(new_n873_), .A3(new_n588_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n902_), .A2(new_n903_), .A3(G134gat), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n882_), .A2(new_n885_), .A3(G134gat), .A4(new_n653_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n902_), .B2(G134gat), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(G1343gat));
  NOR4_X1   g706(.A1(new_n666_), .A2(new_n693_), .A3(new_n334_), .A4(new_n684_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n879_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n658_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n371_), .ZN(G1344gat));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n758_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n372_), .ZN(G1345gat));
  AND2_X1   g712(.A1(new_n879_), .A2(new_n908_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(new_n915_), .A3(new_n529_), .ZN(new_n916_));
  OAI21_X1  g715(.A(KEYINPUT125), .B1(new_n909_), .B2(new_n530_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT61), .B(G155gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1346gat));
  OR3_X1    g719(.A1(new_n909_), .A2(G162gat), .A3(new_n588_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G162gat), .B1(new_n909_), .B2(new_n704_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1347gat));
  AOI21_X1  g722(.A(new_n870_), .B1(new_n319_), .B2(new_n333_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n665_), .A2(new_n446_), .A3(new_n362_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n924_), .A2(new_n646_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n926_), .A2(new_n927_), .A3(G169gat), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n209_), .A2(new_n210_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n926_), .A2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n927_), .B1(new_n926_), .B2(G169gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n928_), .B1(new_n930_), .B2(new_n931_), .ZN(G1348gat));
  NAND2_X1  g731(.A1(new_n924_), .A2(new_n925_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n758_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n277_), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n933_), .A2(new_n530_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n268_), .A2(new_n271_), .B1(new_n937_), .B2(new_n264_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n937_), .A2(G183gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n936_), .B2(new_n940_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n933_), .B2(new_n704_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n589_), .A2(new_n281_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n933_), .B2(new_n943_), .ZN(G1351gat));
  AND2_X1   g743(.A1(new_n448_), .A2(new_n362_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n924_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n658_), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT127), .B(G197gat), .Z(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1352gat));
  NAND3_X1  g748(.A1(new_n924_), .A2(new_n656_), .A3(new_n945_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n924_), .A2(new_n529_), .A3(new_n945_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  AND2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n952_), .A2(new_n953_), .A3(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n952_), .B2(new_n953_), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n946_), .B2(new_n704_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n589_), .A2(new_n232_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n946_), .B2(new_n958_), .ZN(G1355gat));
endmodule


