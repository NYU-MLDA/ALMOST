//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT92), .B1(new_n203_), .B2(G197gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT92), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(new_n206_), .A3(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n203_), .A2(G197gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(new_n203_), .B2(G197gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n206_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(new_n209_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT21), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n204_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n211_), .A2(new_n208_), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n212_), .A2(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT25), .B(G183gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT26), .B(G190gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n228_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT98), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(KEYINPUT22), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT22), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G169gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n241_), .A3(new_n230_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n232_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT97), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(KEYINPUT97), .A3(new_n232_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n238_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n242_), .A2(KEYINPUT97), .A3(new_n232_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT97), .B1(new_n242_), .B2(new_n232_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n238_), .B(new_n252_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n220_), .B(new_n237_), .C1(new_n253_), .C2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT100), .ZN(new_n259_));
  INV_X1    g058(.A(new_n237_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n252_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT98), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n262_), .B2(new_n256_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT100), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n220_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT20), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n251_), .B1(new_n243_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n242_), .A2(KEYINPUT84), .A3(new_n232_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n231_), .A2(new_n232_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n274_), .B2(KEYINPUT24), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n271_), .A2(new_n272_), .B1(new_n228_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT99), .B1(new_n276_), .B2(new_n220_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT99), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n217_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n219_), .A2(new_n218_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n272_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT84), .B1(new_n242_), .B2(new_n232_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n251_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n275_), .A2(new_n228_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n278_), .B(new_n281_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n269_), .B1(new_n277_), .B2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n259_), .A2(new_n265_), .A3(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G8gat), .B(G36gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT18), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G64gat), .B(G92gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT20), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n276_), .B2(new_n220_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(new_n263_), .B2(new_n220_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n267_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(new_n292_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT106), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT106), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n288_), .A2(new_n296_), .A3(new_n299_), .A4(new_n292_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n268_), .B(new_n294_), .C1(new_n263_), .C2(new_n220_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n261_), .A2(new_n237_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT20), .B1(new_n303_), .B2(new_n281_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n277_), .B2(new_n286_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n302_), .B1(new_n305_), .B2(new_n268_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n292_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n301_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n298_), .A2(new_n300_), .A3(new_n308_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n288_), .A2(new_n292_), .A3(new_n296_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n292_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n301_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT1), .ZN(new_n318_));
  INV_X1    g117(.A(G155gat), .ZN(new_n319_));
  INV_X1    g118(.A(G162gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n316_), .B(new_n318_), .C1(new_n323_), .C2(KEYINPUT1), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328_));
  INV_X1    g127(.A(G141gat), .ZN(new_n329_));
  INV_X1    g128(.A(G148gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  AND4_X1   g132(.A1(new_n327_), .A2(new_n331_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT87), .B1(new_n317_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n321_), .A2(new_n337_), .A3(new_n322_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n324_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n343_));
  INV_X1    g142(.A(G134gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G127gat), .ZN(new_n345_));
  INV_X1    g144(.A(G127gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G134gat), .ZN(new_n347_));
  INV_X1    g146(.A(G120gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G113gat), .ZN(new_n349_));
  INV_X1    g148(.A(G113gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G120gat), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n345_), .A2(new_n347_), .A3(new_n349_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n345_), .A2(new_n347_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n343_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n345_), .A2(new_n347_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n349_), .A2(new_n351_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n352_), .A3(KEYINPUT86), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n331_), .A2(new_n327_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(KEYINPUT88), .A3(new_n324_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n342_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n324_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT101), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n364_), .A2(new_n366_), .A3(KEYINPUT101), .A4(KEYINPUT4), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT102), .B(KEYINPUT4), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n342_), .A2(new_n360_), .A3(new_n363_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n364_), .A2(new_n366_), .A3(new_n374_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G85gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT0), .B(G57gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n383_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n376_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n379_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT105), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n386_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395_));
  INV_X1    g194(.A(new_n363_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT88), .B1(new_n362_), .B2(new_n324_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT28), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n342_), .A2(new_n363_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT28), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n395_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G22gat), .B(G50gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT89), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n404_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n281_), .B1(new_n365_), .B2(new_n395_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(KEYINPUT94), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT94), .ZN(new_n416_));
  AOI22_X1  g215(.A1(KEYINPUT29), .A2(new_n340_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n413_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n413_), .B(KEYINPUT90), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n220_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n342_), .A2(KEYINPUT29), .A3(new_n363_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n419_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(KEYINPUT95), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n427_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n419_), .B(new_n429_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT95), .B1(new_n426_), .B2(new_n427_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n411_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n426_), .A2(new_n427_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(new_n430_), .A3(new_n404_), .A4(new_n408_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n313_), .A2(new_n394_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT107), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n313_), .A2(new_n394_), .A3(new_n436_), .A4(KEYINPUT107), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT103), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n373_), .A2(new_n374_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n371_), .A2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n364_), .A2(new_n366_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n383_), .B1(new_n444_), .B2(new_n375_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n384_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n378_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n388_), .B2(new_n384_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n288_), .A2(new_n296_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n307_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n297_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n441_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n386_), .A2(new_n390_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n306_), .A2(KEYINPUT32), .A3(new_n292_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n292_), .A2(KEYINPUT32), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT104), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n456_), .B(new_n457_), .C1(new_n452_), .C2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n310_), .A2(new_n311_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n378_), .A2(new_n448_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT103), .A4(new_n450_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n455_), .A2(new_n460_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n436_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n439_), .A2(new_n440_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT85), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT30), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(new_n276_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n472_), .B(G71gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n471_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n360_), .B(KEYINPUT31), .ZN(new_n475_));
  INV_X1    g274(.A(G99gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n477_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n467_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT108), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT109), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n313_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n313_), .A2(new_n483_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n394_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(new_n480_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n465_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT108), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n467_), .A2(new_n490_), .A3(new_n480_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n482_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G190gat), .B(G218gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G134gat), .B(G162gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(KEYINPUT36), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT34), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(KEYINPUT67), .A3(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(KEYINPUT67), .B2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT6), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(new_n515_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n513_), .B(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n511_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n520_), .B1(new_n524_), .B2(new_n515_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n518_), .A2(KEYINPUT64), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT64), .B1(new_n518_), .B2(new_n526_), .ZN(new_n528_));
  OAI221_X1 g327(.A(new_n517_), .B1(new_n526_), .B2(new_n518_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT65), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT10), .B(G99gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n513_), .B1(G106gat), .B2(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT75), .ZN(new_n535_));
  XOR2_X1   g334(.A(G29gat), .B(G36gat), .Z(new_n536_));
  XOR2_X1   g335(.A(G43gat), .B(G50gat), .Z(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n534_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n538_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n525_), .A2(new_n542_), .A3(new_n533_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n500_), .A2(new_n501_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n535_), .B1(new_n534_), .B2(new_n540_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n502_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n543_), .A2(new_n544_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n502_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .A4(new_n541_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT76), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n497_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n547_), .A2(new_n551_), .A3(KEYINPUT76), .A4(new_n496_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(KEYINPUT36), .A3(new_n495_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT110), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(KEYINPUT110), .A3(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT83), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565_));
  INV_X1    g364(.A(G8gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G1gat), .B(G8gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n538_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n538_), .A2(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(KEYINPUT79), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT79), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n538_), .A2(new_n576_), .A3(new_n570_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT80), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n540_), .A2(new_n570_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n574_), .A3(new_n571_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT81), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT81), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n580_), .A2(new_n583_), .A3(new_n574_), .A4(new_n571_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n579_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n564_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n579_), .A2(new_n585_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n588_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n590_), .A3(new_n564_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n594_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n595_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n591_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G57gat), .B(G64gat), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT11), .ZN(new_n605_));
  XOR2_X1   g404(.A(G71gat), .B(G78gat), .Z(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n604_), .A2(KEYINPUT11), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n606_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT70), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n525_), .A3(new_n533_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n525_), .B2(new_n533_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n603_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT5), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n610_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n534_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n623_), .B(new_n612_), .C1(new_n614_), .C2(KEYINPUT12), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n615_), .B(new_n619_), .C1(new_n624_), .C2(new_n603_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT72), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n534_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n620_), .B1(new_n628_), .B2(new_n611_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n629_), .A2(new_n602_), .A3(new_n612_), .A4(new_n623_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(KEYINPUT72), .A3(new_n615_), .A4(new_n619_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT73), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n615_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n619_), .B(KEYINPUT71), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n632_), .A2(new_n633_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n633_), .B1(new_n632_), .B2(new_n637_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n601_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(KEYINPUT13), .A3(new_n638_), .ZN(new_n643_));
  XOR2_X1   g442(.A(G127gat), .B(G155gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT17), .ZN(new_n649_));
  INV_X1    g448(.A(new_n611_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n570_), .B(new_n651_), .Z(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n653_), .A2(new_n610_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n610_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n656_), .A2(KEYINPUT17), .A3(new_n648_), .A4(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AND4_X1   g459(.A1(new_n600_), .A2(new_n641_), .A3(new_n643_), .A4(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n492_), .A2(new_n563_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n202_), .B1(new_n663_), .B2(new_n487_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n492_), .A2(new_n600_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n641_), .A2(new_n643_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n558_), .B(KEYINPUT37), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n659_), .B(KEYINPUT78), .Z(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(new_n666_), .A3(new_n670_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n671_), .A2(G1gat), .A3(new_n394_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT38), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n664_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n673_), .B2(new_n672_), .ZN(G1324gat));
  INV_X1    g474(.A(new_n486_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n492_), .A2(new_n676_), .A3(new_n563_), .A4(new_n661_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(G8gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n677_), .B2(G8gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(new_n566_), .ZN(new_n682_));
  OAI22_X1  g481(.A1(new_n680_), .A2(new_n681_), .B1(new_n671_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT111), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI221_X1 g484(.A(KEYINPUT111), .B1(new_n671_), .B2(new_n682_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1325gat));
  INV_X1    g489(.A(new_n480_), .ZN(new_n691_));
  INV_X1    g490(.A(G15gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n671_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n663_), .B2(new_n691_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT113), .B(KEYINPUT41), .Z(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(new_n695_), .B2(new_n696_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n662_), .B2(new_n465_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n465_), .A2(G22gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n671_), .B2(new_n701_), .ZN(G1327gat));
  NAND2_X1  g501(.A1(new_n641_), .A2(new_n643_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n563_), .A2(new_n703_), .A3(new_n668_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n665_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n487_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n491_), .A2(new_n489_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n490_), .B1(new_n467_), .B2(new_n480_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n667_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT114), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n558_), .A2(KEYINPUT37), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT37), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT43), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n710_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n492_), .A2(new_n667_), .A3(new_n716_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n600_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n703_), .A2(new_n721_), .A3(new_n668_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT44), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724_));
  INV_X1    g523(.A(new_n722_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n724_), .B(new_n725_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n723_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n487_), .A2(G29gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n707_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n727_), .B2(new_n676_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT115), .B(KEYINPUT45), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n486_), .A2(G36gat), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  OR3_X1    g534(.A1(new_n705_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n733_), .B1(new_n705_), .B2(new_n735_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n730_), .B1(new_n732_), .B2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n736_), .A2(new_n737_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n723_), .A2(new_n726_), .A3(new_n486_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n740_), .B(KEYINPUT46), .C1(new_n741_), .C2(new_n731_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1329gat));
  NAND2_X1  g542(.A1(new_n691_), .A2(G43gat), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n723_), .A2(new_n726_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G43gat), .B1(new_n706_), .B2(new_n691_), .ZN(new_n746_));
  OR3_X1    g545(.A1(new_n745_), .A2(KEYINPUT47), .A3(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT47), .B1(new_n745_), .B2(new_n746_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1330gat));
  OR3_X1    g548(.A1(new_n705_), .A2(G50gat), .A3(new_n465_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n727_), .A2(KEYINPUT116), .A3(new_n436_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT116), .B1(new_n727_), .B2(new_n436_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1331gat));
  NOR3_X1   g553(.A1(new_n666_), .A2(new_n600_), .A3(new_n669_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n492_), .A3(new_n563_), .ZN(new_n756_));
  INV_X1    g555(.A(G57gat), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n394_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n492_), .A2(new_n721_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n666_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT117), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT117), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n487_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n758_), .B1(new_n765_), .B2(new_n757_), .ZN(G1332gat));
  OAI21_X1  g565(.A(G64gat), .B1(new_n756_), .B2(new_n486_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT48), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n486_), .A2(G64gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n761_), .B2(new_n769_), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n756_), .B2(new_n480_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT49), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n480_), .A2(G71gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n761_), .B2(new_n773_), .ZN(G1334gat));
  OAI21_X1  g573(.A(G78gat), .B1(new_n756_), .B2(new_n465_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT50), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n465_), .A2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n761_), .B2(new_n777_), .ZN(G1335gat));
  NOR3_X1   g577(.A1(new_n666_), .A2(new_n600_), .A3(new_n668_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n720_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780_), .B2(new_n394_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n759_), .A2(new_n703_), .A3(new_n669_), .A4(new_n562_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n394_), .A2(G85gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n780_), .B2(new_n486_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n486_), .A2(G92gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n782_), .B2(new_n786_), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n780_), .B2(new_n480_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n480_), .A2(new_n531_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n782_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n790_), .B(new_n792_), .ZN(G1338gat));
  OR3_X1    g592(.A1(new_n782_), .A2(G106gat), .A3(new_n465_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n720_), .A2(new_n436_), .A3(new_n779_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(G106gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n795_), .B2(G106gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n794_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  AND3_X1   g602(.A1(new_n596_), .A2(new_n599_), .A3(new_n632_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n624_), .A2(new_n603_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n630_), .A2(new_n805_), .A3(KEYINPUT55), .ZN(new_n806_));
  OR3_X1    g605(.A1(new_n624_), .A2(KEYINPUT55), .A3(new_n603_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n635_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n807_), .A3(KEYINPUT120), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n811_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n804_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n580_), .A2(new_n575_), .A3(new_n571_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n573_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n594_), .A3(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n589_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n562_), .B1(new_n814_), .B2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n632_), .A2(new_n818_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT58), .B(new_n821_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n667_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n808_), .A2(new_n809_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n636_), .A3(new_n811_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n811_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT58), .B1(new_n829_), .B2(new_n821_), .ZN(new_n830_));
  OAI22_X1  g629(.A1(new_n820_), .A2(KEYINPUT57), .B1(new_n823_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n814_), .A2(new_n819_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT57), .A3(new_n563_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n659_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n836_));
  NOR2_X1   g635(.A1(new_n712_), .A2(new_n714_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n666_), .A2(new_n837_), .A3(new_n668_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n838_), .B2(new_n600_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT54), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n670_), .A2(new_n666_), .A3(new_n721_), .A4(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n835_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n486_), .A2(new_n691_), .A3(new_n487_), .A4(new_n465_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(new_n350_), .A3(new_n600_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(KEYINPUT59), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n669_), .B1(new_n831_), .B2(new_n834_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n843_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n846_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n850_), .A2(new_n600_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n849_), .B1(new_n855_), .B2(new_n350_), .ZN(G1340gat));
  OAI21_X1  g655(.A(new_n348_), .B1(new_n666_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n848_), .B(new_n857_), .C1(KEYINPUT60), .C2(new_n348_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n850_), .A2(new_n703_), .A3(new_n854_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n348_), .ZN(G1341gat));
  NAND3_X1  g659(.A1(new_n848_), .A2(new_n346_), .A3(new_n668_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n850_), .A2(new_n660_), .A3(new_n854_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n346_), .ZN(G1342gat));
  NAND3_X1  g662(.A1(new_n848_), .A2(new_n344_), .A3(new_n562_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n850_), .A2(new_n667_), .A3(new_n854_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n344_), .ZN(G1343gat));
  AOI21_X1  g665(.A(new_n691_), .B1(new_n835_), .B2(new_n843_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n676_), .A2(new_n394_), .A3(new_n465_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n721_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n329_), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n666_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT121), .B(G148gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1345gat));
  NOR2_X1   g673(.A1(new_n869_), .A2(new_n669_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n875_), .B(new_n877_), .ZN(G1346gat));
  AND2_X1   g677(.A1(new_n867_), .A2(new_n868_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G162gat), .B1(new_n879_), .B2(new_n562_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n667_), .A2(G162gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT122), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n879_), .B2(new_n882_), .ZN(G1347gat));
  NAND3_X1  g682(.A1(new_n676_), .A2(new_n465_), .A3(new_n488_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n851_), .B2(new_n843_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n229_), .B1(new_n885_), .B2(new_n600_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n885_), .A2(new_n239_), .A3(new_n241_), .A4(new_n600_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(G1348gat));
  AOI21_X1  g689(.A(new_n884_), .B1(new_n835_), .B2(new_n843_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n666_), .A2(new_n230_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT124), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n895_), .A3(new_n892_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898_));
  INV_X1    g697(.A(new_n885_), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n898_), .B(new_n230_), .C1(new_n899_), .C2(new_n666_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n666_), .B(new_n884_), .C1(new_n851_), .C2(new_n843_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT123), .B1(new_n901_), .B2(G176gat), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n897_), .A2(new_n900_), .A3(new_n902_), .ZN(G1349gat));
  AOI21_X1  g702(.A(G183gat), .B1(new_n891_), .B2(new_n668_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n659_), .A2(new_n226_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n885_), .B2(new_n905_), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n899_), .B2(new_n837_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n885_), .A2(new_n227_), .A3(new_n562_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1351gat));
  NOR2_X1   g708(.A1(new_n487_), .A2(new_n465_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n676_), .A2(new_n910_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n691_), .B(new_n911_), .C1(new_n835_), .C2(new_n843_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n600_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n703_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g715(.A(new_n659_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n912_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n919_), .A2(KEYINPUT125), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n919_), .B(KEYINPUT125), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n918_), .B2(new_n922_), .ZN(G1354gat));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n924_));
  AOI21_X1  g723(.A(G218gat), .B1(new_n912_), .B2(new_n562_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n911_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n667_), .A2(G218gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT126), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n867_), .A2(new_n926_), .A3(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n924_), .B1(new_n925_), .B2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n912_), .A2(new_n928_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n867_), .A2(new_n562_), .A3(new_n926_), .ZN(new_n932_));
  OAI211_X1 g731(.A(KEYINPUT127), .B(new_n931_), .C1(new_n932_), .C2(G218gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n930_), .A2(new_n933_), .ZN(G1355gat));
endmodule


