//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n815_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT19), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT20), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n205_), .B1(G183gat), .B2(G190gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT81), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT81), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n209_), .A2(new_n205_), .A3(G183gat), .A4(G190gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n206_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n212_), .A2(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n218_));
  OR2_X1    g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n211_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT95), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n218_), .A2(KEYINPUT95), .A3(new_n222_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n219_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n206_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n207_), .A2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n205_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n232_), .A2(new_n234_), .B1(G169gat), .B2(G176gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n221_), .A2(new_n227_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G211gat), .B(G218gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT21), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G197gat), .B(G204gat), .Z(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n240_), .A2(KEYINPUT21), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n245_), .A2(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n246_), .B2(new_n243_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n204_), .B1(new_n239_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n208_), .A2(new_n210_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n228_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n234_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT82), .B1(new_n211_), .B2(new_n233_), .ZN(new_n253_));
  AOI21_X1  g052(.A(G176gat), .B1(KEYINPUT80), .B2(KEYINPUT22), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G169gat), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT78), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n216_), .A2(KEYINPUT77), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(G190gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n222_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n257_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  AOI211_X1 g065(.A(KEYINPUT78), .B(new_n266_), .C1(new_n258_), .C2(new_n262_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n232_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n256_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n203_), .B(new_n248_), .C1(new_n271_), .C2(new_n247_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT96), .ZN(new_n273_));
  INV_X1    g072(.A(new_n262_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n261_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n264_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT78), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n263_), .A2(new_n257_), .A3(new_n264_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n270_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n247_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n239_), .A2(new_n247_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT20), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n203_), .B(KEYINPUT93), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n280_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n247_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT96), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n203_), .A4(new_n248_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n273_), .A2(new_n285_), .A3(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT98), .ZN(new_n293_));
  XOR2_X1   g092(.A(G64gat), .B(G92gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n298_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n273_), .A2(new_n285_), .A3(new_n297_), .A4(new_n290_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(KEYINPUT99), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302_));
  INV_X1    g101(.A(new_n291_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT99), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(new_n297_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT102), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n301_), .A2(new_n305_), .A3(KEYINPUT102), .A4(new_n302_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G113gat), .B(G120gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT85), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G127gat), .B(G134gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT84), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n316_), .B(KEYINPUT84), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n314_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n320_), .A3(KEYINPUT86), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n319_), .A2(KEYINPUT86), .A3(new_n314_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(KEYINPUT89), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT88), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT89), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n326_), .B(new_n328_), .Z(new_n329_));
  NAND2_X1  g128(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n330_));
  OR2_X1    g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n330_), .A3(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n339_), .B2(new_n335_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n325_), .A3(new_n331_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n323_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n342_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n318_), .A2(new_n320_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n349_), .A2(KEYINPUT4), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT4), .B1(new_n323_), .B2(new_n343_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n312_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n344_), .A2(new_n311_), .A3(new_n348_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n351_), .B1(new_n349_), .B2(KEYINPUT4), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n353_), .B(new_n358_), .C1(new_n361_), .C2(new_n311_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n287_), .B1(new_n346_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G106gat), .ZN(new_n366_));
  INV_X1    g165(.A(G106gat), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n367_), .B(new_n287_), .C1(new_n346_), .C2(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G78gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT92), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n366_), .A2(new_n372_), .A3(new_n368_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n374_), .A2(KEYINPUT90), .A3(new_n376_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n375_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n346_), .A2(new_n364_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT28), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(KEYINPUT28), .ZN(new_n383_));
  OAI21_X1  g182(.A(G22gat), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  INV_X1    g184(.A(G22gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n381_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n387_), .A3(G50gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(G50gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n379_), .A2(new_n388_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n388_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n363_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n288_), .A2(new_n248_), .ZN(new_n396_));
  OAI22_X1  g195(.A1(new_n396_), .A2(new_n203_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n298_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n300_), .A3(KEYINPUT27), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n310_), .A2(new_n395_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT103), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n301_), .A2(new_n305_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n352_), .A2(new_n403_), .A3(new_n353_), .A4(new_n358_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n362_), .A2(KEYINPUT33), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n344_), .A2(new_n312_), .A3(new_n348_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n407_), .B(new_n359_), .C1(new_n361_), .C2(new_n312_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n402_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT100), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n402_), .A2(new_n406_), .A3(new_n411_), .A4(new_n408_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n297_), .A2(KEYINPUT32), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n397_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT101), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n415_), .B(new_n363_), .C1(new_n291_), .C2(new_n413_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n410_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n392_), .A2(new_n394_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n399_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT103), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n395_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n401_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n323_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G71gat), .B(G99gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT31), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G15gat), .B(G43gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n286_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n429_), .B(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(new_n363_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n422_), .A2(new_n419_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT104), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n422_), .A2(KEYINPUT104), .A3(new_n419_), .A4(new_n436_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n425_), .A2(new_n435_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G22gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G1gat), .A2(G8gat), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n443_), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT74), .B1(new_n443_), .B2(KEYINPUT14), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n442_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G8gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G231gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G57gat), .B(G64gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT11), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G71gat), .B(G78gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n452_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n451_), .A2(KEYINPUT11), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n454_), .B1(new_n457_), .B2(new_n453_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n450_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G127gat), .B(G155gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G211gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT16), .B(G183gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n462_), .B(new_n463_), .Z(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(KEYINPUT17), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n464_), .A2(new_n466_), .A3(KEYINPUT17), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n465_), .B(new_n467_), .Z(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G232gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT34), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT35), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT69), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  XOR2_X1   g273(.A(G85gat), .B(G92gat), .Z(new_n475_));
  NAND2_X1  g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT6), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT65), .ZN(new_n478_));
  NOR2_X1   g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n482_), .B2(new_n480_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n474_), .B(new_n475_), .C1(new_n478_), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n477_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n475_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT8), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT9), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n475_), .B2(new_n492_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT64), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(KEYINPUT64), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n478_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT10), .B(G99gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n490_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G29gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  XOR2_X1   g303(.A(new_n504_), .B(KEYINPUT15), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  OAI22_X1  g305(.A1(new_n506_), .A2(KEYINPUT70), .B1(KEYINPUT35), .B2(new_n471_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(KEYINPUT70), .B2(new_n506_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n501_), .A2(new_n504_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT71), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n473_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G190gat), .B(G218gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G162gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT72), .B(G134gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n506_), .A2(new_n473_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n471_), .A2(KEYINPUT35), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n510_), .A2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n512_), .A2(new_n513_), .A3(new_n517_), .A4(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n513_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n517_), .A2(new_n513_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n521_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n523_), .B(new_n524_), .C1(new_n525_), .C2(new_n511_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT37), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n526_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT73), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n441_), .A2(new_n469_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n505_), .A2(new_n448_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT75), .B1(new_n448_), .B2(new_n504_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n537_), .B(new_n538_), .C1(new_n539_), .C2(new_n535_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n448_), .B(new_n504_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(G229gat), .A3(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT76), .B(G169gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G197gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n540_), .A2(new_n542_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT67), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n501_), .A2(new_n555_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n489_), .A2(new_n486_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n554_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n558_), .A3(new_n458_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n501_), .A2(new_n466_), .A3(KEYINPUT12), .A4(new_n459_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n553_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n557_), .B(new_n459_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n553_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT5), .B(G176gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G204gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G120gat), .B(G148gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n562_), .A2(new_n564_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT13), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n573_), .A2(new_n574_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT68), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n534_), .A2(new_n551_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(G1gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n363_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT105), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n425_), .A2(new_n435_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n439_), .A2(new_n440_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n468_), .A3(new_n530_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n551_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n578_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n363_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n586_), .A2(new_n587_), .A3(new_n597_), .ZN(G1324gat));
  INV_X1    g397(.A(G8gat), .ZN(new_n599_));
  INV_X1    g398(.A(new_n422_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n581_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n594_), .A2(new_n600_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(G8gat), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(KEYINPUT39), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(KEYINPUT39), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n601_), .B(new_n607_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1325gat));
  INV_X1    g410(.A(G15gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n435_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n594_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT41), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n581_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1326gat));
  AOI21_X1  g416(.A(new_n386_), .B1(new_n594_), .B2(new_n418_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT42), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n581_), .A2(new_n386_), .A3(new_n418_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1327gat));
  INV_X1    g420(.A(new_n533_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT43), .B1(new_n441_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT43), .ZN(new_n624_));
  AND4_X1   g423(.A1(new_n423_), .A2(new_n310_), .A3(new_n395_), .A4(new_n399_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n423_), .B1(new_n422_), .B2(new_n395_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n613_), .B1(new_n627_), .B2(new_n420_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n589_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n624_), .B(new_n533_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n593_), .A2(new_n592_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n469_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT44), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  AOI211_X1 g435(.A(new_n636_), .B(new_n633_), .C1(new_n623_), .C2(new_n630_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n363_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT107), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT107), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n641_), .A3(new_n363_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(G29gat), .A3(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n441_), .A2(new_n530_), .A3(new_n633_), .ZN(new_n644_));
  INV_X1    g443(.A(G29gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n363_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(G1328gat));
  INV_X1    g446(.A(G36gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n648_), .A3(new_n600_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT109), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n644_), .A2(KEYINPUT109), .A3(new_n648_), .A4(new_n600_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n635_), .A2(new_n637_), .A3(new_n422_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n655_), .B(KEYINPUT46), .C1(new_n648_), .C2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  INV_X1    g457(.A(new_n654_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n653_), .B(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n656_), .A2(new_n648_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n662_), .ZN(G1329gat));
  NAND2_X1  g462(.A1(new_n644_), .A2(new_n613_), .ZN(new_n664_));
  INV_X1    g463(.A(G43gat), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n435_), .A2(new_n665_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n638_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n668_), .ZN(new_n670_));
  NOR4_X1   g469(.A1(new_n635_), .A2(new_n637_), .A3(KEYINPUT110), .A4(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT47), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT47), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n674_), .B(new_n666_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1330gat));
  NOR3_X1   g475(.A1(new_n635_), .A2(new_n637_), .A3(new_n419_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n677_), .A2(KEYINPUT111), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(KEYINPUT111), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(G50gat), .A3(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n644_), .A2(new_n390_), .A3(new_n418_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1331gat));
  AND3_X1   g481(.A1(new_n534_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n363_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n579_), .A2(new_n592_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n591_), .A2(new_n596_), .A3(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(G57gat), .B2(new_n686_), .ZN(G1332gat));
  INV_X1    g486(.A(G64gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n591_), .A2(new_n685_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n600_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT48), .Z(new_n691_));
  NAND3_X1  g490(.A1(new_n683_), .A2(new_n688_), .A3(new_n600_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1333gat));
  INV_X1    g492(.A(G71gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n689_), .B2(new_n613_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT49), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n683_), .A2(new_n694_), .A3(new_n613_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1334gat));
  AOI21_X1  g497(.A(new_n371_), .B1(new_n689_), .B2(new_n418_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT50), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n683_), .A2(new_n371_), .A3(new_n418_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1335gat));
  NAND3_X1  g501(.A1(new_n590_), .A2(new_n469_), .A3(new_n527_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n685_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G85gat), .B1(new_n704_), .B2(new_n363_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n578_), .A2(new_n551_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n631_), .A2(new_n469_), .A3(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n363_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n705_), .B1(new_n708_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g508(.A(new_n704_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n710_), .A2(G92gat), .A3(new_n422_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n600_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(G92gat), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT112), .ZN(G1337gat));
  NOR3_X1   g513(.A1(new_n710_), .A2(new_n498_), .A3(new_n435_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n707_), .A2(new_n613_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(G99gat), .B2(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g517(.A1(new_n704_), .A2(new_n367_), .A3(new_n418_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n631_), .A2(new_n469_), .A3(new_n418_), .A4(new_n706_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(G106gat), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n720_), .B2(G106gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g524(.A1(new_n528_), .A2(new_n532_), .A3(new_n592_), .A4(new_n468_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n726_), .A2(new_n593_), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n726_), .B2(new_n593_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT56), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n559_), .A2(new_n560_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n552_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n562_), .A2(KEYINPUT55), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT55), .B(new_n553_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n734_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n732_), .B1(new_n738_), .B2(new_n571_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT116), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n561_), .A2(new_n741_), .ZN(new_n742_));
  OAI22_X1  g541(.A1(new_n742_), .A2(new_n736_), .B1(new_n552_), .B2(new_n733_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(KEYINPUT56), .A3(new_n569_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n740_), .A3(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n743_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n569_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(new_n572_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n541_), .A2(new_n538_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n537_), .B1(new_n539_), .B2(new_n535_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n547_), .B(new_n748_), .C1(new_n749_), .C2(new_n538_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n550_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n747_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT58), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n745_), .A2(new_n747_), .A3(KEYINPUT58), .A4(new_n751_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n533_), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n739_), .A2(new_n744_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n572_), .A2(new_n551_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT115), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n759_), .A2(new_n761_), .B1(new_n573_), .B2(new_n751_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n762_), .B2(new_n527_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(new_n761_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n573_), .A2(new_n751_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(KEYINPUT57), .A3(new_n530_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n756_), .A2(new_n757_), .A3(new_n763_), .A4(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n469_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n767_), .A2(new_n763_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n757_), .B1(new_n770_), .B2(new_n756_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n731_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n422_), .A2(new_n363_), .A3(new_n613_), .A4(new_n419_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT118), .Z(new_n774_));
  AND2_X1   g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G113gat), .B1(new_n775_), .B2(new_n551_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n729_), .A2(new_n730_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n468_), .B1(new_n770_), .B2(new_n756_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n774_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n772_), .A2(new_n774_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(KEYINPUT59), .B2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(new_n551_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n776_), .B1(new_n785_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n784_), .A2(new_n787_), .A3(new_n579_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n784_), .B2(new_n579_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G120gat), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT60), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n578_), .B2(G120gat), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n775_), .B(new_n792_), .C1(new_n791_), .C2(G120gat), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1341gat));
  AOI21_X1  g593(.A(G127gat), .B1(new_n775_), .B2(new_n468_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n784_), .A2(G127gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n468_), .ZN(G1342gat));
  AOI21_X1  g596(.A(G134gat), .B1(new_n775_), .B2(new_n527_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT120), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n784_), .A2(G134gat), .A3(new_n533_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1343gat));
  NOR2_X1   g600(.A1(new_n600_), .A2(new_n613_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n772_), .A2(new_n363_), .A3(new_n418_), .A4(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n756_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n767_), .A2(new_n763_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT117), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n469_), .A3(new_n768_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n419_), .B1(new_n809_), .B2(new_n731_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n810_), .A2(KEYINPUT121), .A3(new_n363_), .A4(new_n802_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n805_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n551_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n579_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n468_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT61), .B(G155gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n817_), .B(new_n818_), .ZN(G1346gat));
  NAND2_X1  g618(.A1(new_n533_), .A2(G162gat), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT123), .Z(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n805_), .B2(new_n811_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n812_), .A2(new_n527_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  INV_X1    g623(.A(G162gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n530_), .B1(new_n805_), .B2(new_n811_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT122), .B1(new_n827_), .B2(G162gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n822_), .B1(new_n826_), .B2(new_n828_), .ZN(G1347gat));
  INV_X1    g628(.A(new_n779_), .ZN(new_n830_));
  NOR4_X1   g629(.A1(new_n422_), .A2(new_n363_), .A3(new_n435_), .A4(new_n418_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n551_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(G169gat), .A3(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n551_), .A2(new_n236_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT125), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n839_), .A2(KEYINPUT125), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n833_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n837_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n834_), .A2(G169gat), .A3(new_n843_), .A4(new_n835_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n838_), .A2(new_n842_), .A3(new_n844_), .ZN(G1348gat));
  NAND4_X1  g644(.A1(new_n772_), .A2(G176gat), .A3(new_n579_), .A4(new_n831_), .ZN(new_n846_));
  XOR2_X1   g645(.A(new_n846_), .B(KEYINPUT126), .Z(new_n847_));
  AOI21_X1  g646(.A(G176gat), .B1(new_n833_), .B2(new_n593_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1349gat));
  NOR2_X1   g648(.A1(new_n832_), .A2(new_n469_), .ZN(new_n850_));
  MUX2_X1   g649(.A(G183gat), .B(new_n259_), .S(new_n850_), .Z(G1350gat));
  OAI21_X1  g650(.A(G190gat), .B1(new_n832_), .B2(new_n622_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n527_), .A2(new_n260_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n832_), .B2(new_n853_), .ZN(G1351gat));
  AOI211_X1 g653(.A(new_n613_), .B(new_n422_), .C1(new_n809_), .C2(new_n731_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n855_), .A2(new_n395_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n551_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n579_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G204gat), .ZN(G1353gat));
  AND3_X1   g659(.A1(new_n855_), .A2(new_n468_), .A3(new_n395_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n861_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT63), .B(G211gat), .Z(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n861_), .B2(new_n863_), .ZN(G1354gat));
  NAND3_X1  g663(.A1(new_n855_), .A2(new_n395_), .A3(new_n533_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G218gat), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT127), .ZN(new_n867_));
  INV_X1    g666(.A(G218gat), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n855_), .A2(new_n868_), .A3(new_n527_), .A4(new_n395_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n866_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n866_), .B2(new_n869_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1355gat));
endmodule


