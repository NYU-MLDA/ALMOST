//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n979_, new_n980_, new_n981_, new_n983_, new_n984_,
    new_n985_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n996_, new_n997_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1004_, new_n1005_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G120gat), .B(G148gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT5), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G176gat), .B(G204gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  XNOR2_X1  g006(.A(G57gat), .B(G64gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G71gat), .B(G78gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT11), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n211_));
  INV_X1    g010(.A(new_n209_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n210_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT12), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220_));
  AND2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  INV_X1    g023(.A(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT67), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n219_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G99gat), .ZN(new_n230_));
  INV_X1    g029(.A(G106gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT65), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT7), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT6), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT6), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(G99gat), .A3(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT7), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n239_), .A2(new_n230_), .A3(new_n231_), .A4(KEYINPUT65), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n229_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT8), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n229_), .A2(new_n244_), .A3(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT10), .B(G99gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(G106gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n226_), .A2(KEYINPUT9), .A3(new_n227_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n227_), .A2(KEYINPUT9), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n238_), .A4(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n215_), .B1(new_n246_), .B2(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n229_), .A2(new_n244_), .A3(new_n241_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n244_), .B1(new_n229_), .B2(new_n241_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n215_), .B(new_n252_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n218_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n252_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n216_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n262_), .B2(new_n217_), .ZN(new_n263_));
  AOI211_X1 g062(.A(KEYINPUT68), .B(KEYINPUT12), .C1(new_n261_), .C2(new_n216_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n258_), .B(new_n259_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n256_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n259_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n265_), .A2(KEYINPUT69), .A3(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT69), .B1(new_n265_), .B2(new_n268_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n203_), .B(new_n207_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n207_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n272_), .A3(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(new_n268_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n265_), .A2(KEYINPUT69), .A3(new_n268_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n203_), .B1(new_n279_), .B2(new_n207_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n202_), .B1(new_n274_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n207_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT70), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n273_), .A4(new_n271_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(KEYINPUT71), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G113gat), .B(G141gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G169gat), .B(G197gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT81), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G8gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT14), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT77), .B(G8gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(G1gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(G15gat), .B(G22gat), .Z(new_n298_));
  NOR3_X1   g097(.A1(new_n297_), .A2(KEYINPUT78), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300_));
  AND2_X1   g099(.A1(KEYINPUT77), .A2(G8gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(KEYINPUT77), .A2(G8gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(G1gat), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT14), .ZN(new_n304_));
  INV_X1    g103(.A(new_n298_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n294_), .B1(new_n299_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT78), .B1(new_n297_), .B2(new_n298_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n305_), .A3(new_n300_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n293_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G43gat), .B(G50gat), .Z(new_n312_));
  INV_X1    g111(.A(G36gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G29gat), .ZN(new_n314_));
  INV_X1    g113(.A(G29gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G36gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n316_), .A3(KEYINPUT73), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT73), .B1(new_n314_), .B2(new_n316_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n312_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n315_), .A2(G36gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n313_), .A2(G29gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G43gat), .B(G50gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n317_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n311_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G229gat), .A2(G233gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n307_), .A2(new_n310_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT15), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n318_), .A2(new_n319_), .A3(new_n312_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n325_), .B1(new_n324_), .B2(new_n317_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n320_), .A2(new_n326_), .A3(KEYINPUT15), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n336_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT80), .B1(new_n311_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n330_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n311_), .A2(new_n327_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n329_), .B1(new_n344_), .B2(new_n328_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n292_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n329_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n311_), .B2(new_n327_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n338_), .B1(new_n331_), .B2(new_n337_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n311_), .A2(new_n340_), .A3(KEYINPUT80), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n328_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n347_), .B1(new_n352_), .B2(new_n343_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n291_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n346_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT71), .B1(new_n281_), .B2(new_n284_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n286_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(G15gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT30), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT31), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT23), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(G183gat), .B2(G190gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(G169gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n365_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT24), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT25), .B(G183gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT26), .B(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n380_), .A2(KEYINPUT82), .A3(KEYINPUT24), .A4(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n383_));
  INV_X1    g182(.A(new_n381_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n379_), .A2(new_n382_), .A3(KEYINPUT83), .A4(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n376_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n379_), .A2(new_n386_), .A3(new_n382_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n371_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G71gat), .B(G99gat), .Z(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT84), .B(G43gat), .Z(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G127gat), .B(G134gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT85), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400_));
  INV_X1    g199(.A(G127gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(G134gat), .ZN(new_n402_));
  INV_X1    g201(.A(G134gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(G127gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n400_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G113gat), .B(G120gat), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n399_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n399_), .B2(new_n405_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n389_), .A2(new_n390_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n376_), .A2(new_n387_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n370_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n395_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n397_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n409_), .B1(new_n397_), .B2(new_n413_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n364_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n363_), .A3(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT19), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G204gat), .ZN(new_n426_));
  OR2_X1    g225(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G197gat), .A2(G204gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G211gat), .B(G218gat), .Z(new_n433_));
  NAND4_X1  g232(.A1(new_n430_), .A2(KEYINPUT21), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n427_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT21), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(G197gat), .B2(G204gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n433_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT88), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n435_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT20), .B1(new_n392_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n373_), .B1(new_n375_), .B2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n381_), .A3(new_n380_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT91), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n379_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n450_), .B2(new_n379_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n448_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n370_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n444_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT88), .B1(new_n439_), .B2(new_n440_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n434_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n425_), .B1(new_n446_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n392_), .A2(new_n445_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n424_), .A3(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G8gat), .B(G36gat), .Z(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n460_), .A2(new_n464_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n460_), .B2(new_n464_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n422_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G141gat), .B(G148gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G155gat), .A2(G162gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G155gat), .A2(G162gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(KEYINPUT1), .B2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(KEYINPUT1), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT3), .ZN(new_n481_));
  INV_X1    g280(.A(G141gat), .ZN(new_n482_));
  INV_X1    g281(.A(G148gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G141gat), .A2(G148gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT2), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(new_n487_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G155gat), .B(G162gat), .Z(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(KEYINPUT86), .A3(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n480_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n458_), .B1(new_n474_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n497_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G78gat), .B(G106gat), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n490_), .A2(KEYINPUT86), .A3(new_n491_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT86), .B1(new_n490_), .B2(new_n491_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n478_), .A2(new_n479_), .ZN(new_n504_));
  OAI22_X1  g303(.A1(new_n502_), .A2(new_n503_), .B1(new_n504_), .B2(new_n475_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT28), .B1(new_n505_), .B2(KEYINPUT29), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT28), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n496_), .A2(new_n507_), .A3(new_n474_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G22gat), .B(G50gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT89), .B(new_n501_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n506_), .A2(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n509_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n511_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n500_), .B(new_n514_), .C1(new_n501_), .C2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n497_), .B(new_n498_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n512_), .A2(new_n513_), .A3(new_n501_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n501_), .A2(KEYINPUT89), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n516_), .B2(new_n511_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n519_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n460_), .A2(new_n464_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n469_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n448_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n447_), .A2(new_n384_), .A3(new_n375_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n377_), .A2(new_n378_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT91), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n450_), .A2(new_n451_), .A3(new_n379_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n528_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT95), .B1(new_n533_), .B2(new_n371_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n454_), .A2(new_n535_), .A3(new_n370_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n536_), .A3(new_n445_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n461_), .B1(new_n458_), .B2(new_n412_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n425_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(new_n532_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n371_), .B1(new_n540_), .B2(new_n448_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT20), .B1(new_n541_), .B2(new_n445_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n458_), .A2(new_n412_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n424_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n469_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n527_), .A2(new_n545_), .A3(KEYINPUT27), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G1gat), .B(G29gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G85gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n409_), .A2(new_n505_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n407_), .A2(new_n408_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n496_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n555_), .A3(KEYINPUT4), .ZN(new_n556_));
  OR3_X1    g355(.A1(new_n496_), .A2(new_n554_), .A3(KEYINPUT4), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G225gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n552_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n559_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n565_), .A2(new_n551_), .A3(new_n562_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n473_), .A2(new_n524_), .A3(new_n546_), .A4(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n556_), .A2(new_n559_), .A3(new_n557_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n553_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n552_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT33), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n551_), .B1(new_n565_), .B2(new_n562_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT33), .B(new_n551_), .C1(new_n565_), .C2(new_n562_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n574_), .A2(new_n527_), .A3(new_n470_), .A4(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT32), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n469_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n578_), .B(new_n580_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n542_), .A2(new_n543_), .A3(new_n425_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n541_), .A2(new_n445_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n424_), .B1(new_n538_), .B2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n581_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n579_), .B(new_n585_), .C1(new_n564_), .C2(new_n566_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n524_), .B1(new_n576_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n568_), .B1(new_n587_), .B2(KEYINPUT96), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT96), .ZN(new_n589_));
  AOI211_X1 g388(.A(new_n589_), .B(new_n524_), .C1(new_n576_), .C2(new_n586_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n421_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n567_), .A2(new_n420_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n524_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n592_), .A2(new_n593_), .A3(new_n473_), .A4(new_n546_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT98), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n473_), .A2(new_n546_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n593_), .A4(new_n592_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT79), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n311_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n216_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT16), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n604_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n604_), .A2(new_n610_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n337_), .A2(new_n261_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT34), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n619_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n327_), .B(new_n252_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n615_), .A2(new_n621_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n252_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n622_), .B(new_n623_), .C1(new_n626_), .C2(new_n340_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n620_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT74), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(KEYINPUT36), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n624_), .A2(new_n628_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n632_), .B(KEYINPUT36), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n624_), .A2(new_n628_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT76), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n624_), .A2(new_n628_), .A3(KEYINPUT76), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n636_), .B(KEYINPUT75), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(new_n637_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n634_), .A2(KEYINPUT37), .ZN(new_n644_));
  OAI22_X1  g443(.A1(new_n641_), .A2(KEYINPUT37), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n614_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n358_), .A2(new_n600_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(G1gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n567_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n648_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .A4(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT38), .ZN(new_n654_));
  INV_X1    g453(.A(new_n614_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n641_), .B(KEYINPUT100), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n591_), .B2(new_n599_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n358_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n650_), .B1(new_n658_), .B2(new_n651_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT101), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n654_), .A2(new_n660_), .ZN(G1324gat));
  NOR2_X1   g460(.A1(new_n596_), .A2(new_n296_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n649_), .A2(new_n652_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n596_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n658_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n665_), .A2(new_n666_), .A3(G8gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n665_), .B2(G8gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT40), .B(new_n663_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1325gat));
  AOI21_X1  g472(.A(new_n360_), .B1(new_n658_), .B2(new_n420_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT41), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n649_), .A2(new_n652_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n360_), .A3(new_n420_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n593_), .A2(G22gat), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT103), .Z(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n658_), .A2(new_n524_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(G22gat), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G22gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n600_), .B2(new_n645_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n644_), .B1(new_n637_), .B2(new_n642_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n637_), .A2(new_n638_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n636_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n640_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n634_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT37), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n690_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT43), .B(new_n696_), .C1(new_n591_), .C2(new_n599_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n689_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n358_), .A2(new_n614_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n687_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NOR4_X1   g499(.A1(new_n286_), .A2(new_n357_), .A3(new_n356_), .A4(new_n655_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n701_), .B(KEYINPUT44), .C1(new_n689_), .C2(new_n697_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(new_n651_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n357_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n600_), .A2(new_n705_), .A3(new_n355_), .A4(new_n285_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n656_), .A2(new_n614_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT104), .Z(new_n708_));
  NOR2_X1   g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n651_), .A2(new_n315_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT105), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n704_), .A2(new_n315_), .B1(new_n710_), .B2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(KEYINPUT46), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n700_), .A2(new_n664_), .A3(new_n702_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(G36gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(KEYINPUT46), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n596_), .A2(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n709_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n720_), .ZN(new_n722_));
  NOR4_X1   g521(.A1(new_n706_), .A2(new_n708_), .A3(KEYINPUT106), .A4(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT45), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n708_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n725_), .A2(new_n358_), .A3(new_n600_), .A4(new_n720_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT106), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n709_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n724_), .A2(new_n730_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n717_), .A2(new_n718_), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n718_), .B1(new_n717_), .B2(new_n731_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1329gat));
  NAND4_X1  g533(.A1(new_n700_), .A2(G43gat), .A3(new_n702_), .A4(new_n420_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n710_), .A2(new_n421_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(G43gat), .B2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n709_), .B2(new_n524_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n524_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n703_), .B2(new_n741_), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n705_), .A2(new_n285_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n614_), .A2(new_n355_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n657_), .A3(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n567_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n356_), .A3(new_n600_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n646_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n567_), .A2(G57gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1332gat));
  INV_X1    g550(.A(new_n745_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n664_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(G64gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G64gat), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n596_), .A2(G64gat), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT109), .ZN(new_n758_));
  OAI22_X1  g557(.A1(new_n755_), .A2(new_n756_), .B1(new_n749_), .B2(new_n758_), .ZN(G1333gat));
  NAND2_X1  g558(.A1(new_n752_), .A2(new_n420_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G71gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G71gat), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n421_), .A2(G71gat), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n762_), .A2(new_n763_), .B1(new_n749_), .B2(new_n764_), .ZN(G1334gat));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n752_), .A2(new_n524_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G78gat), .ZN(new_n768_));
  INV_X1    g567(.A(G78gat), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT50), .B(new_n769_), .C1(new_n752_), .C2(new_n524_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n524_), .A2(new_n769_), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n768_), .A2(new_n770_), .B1(new_n749_), .B2(new_n771_), .ZN(G1335gat));
  NAND2_X1  g571(.A1(new_n600_), .A2(new_n645_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT43), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n600_), .A2(new_n688_), .A3(new_n645_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n698_), .A2(KEYINPUT110), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n743_), .A2(new_n356_), .A3(new_n614_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782_), .B2(new_n567_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n748_), .A2(new_n224_), .A3(new_n651_), .A4(new_n725_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1336gat));
  OAI21_X1  g584(.A(G92gat), .B1(new_n782_), .B2(new_n596_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n748_), .A2(new_n225_), .A3(new_n664_), .A4(new_n725_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n782_), .B2(new_n421_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n748_), .A2(new_n247_), .A3(new_n420_), .A4(new_n725_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n792_));
  NAND2_X1  g591(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1338gat));
  NAND4_X1  g594(.A1(new_n748_), .A2(new_n248_), .A3(new_n524_), .A4(new_n725_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n776_), .A2(new_n781_), .A3(new_n524_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n796_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n267_), .B2(KEYINPUT114), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n807_), .B2(new_n267_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n258_), .B(new_n809_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT68), .B1(new_n253_), .B2(KEYINPUT12), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n262_), .A2(new_n260_), .A3(new_n217_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n811_), .A2(new_n812_), .B1(new_n266_), .B2(new_n218_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n808_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n810_), .B(new_n207_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n258_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n808_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n207_), .A4(new_n810_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n328_), .B(new_n347_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n329_), .B1(new_n352_), .B2(new_n343_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n289_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n290_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n273_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n821_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n696_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n826_), .B1(new_n820_), .B2(new_n817_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT117), .B1(new_n831_), .B2(KEYINPUT58), .ZN(new_n832_));
  AND4_X1   g631(.A1(KEYINPUT117), .A2(new_n821_), .A3(KEYINPUT58), .A4(new_n827_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n830_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT118), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n830_), .B(new_n836_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n815_), .A2(KEYINPUT115), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n819_), .A2(new_n841_), .A3(new_n207_), .A4(new_n810_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(new_n816_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n840_), .A2(KEYINPUT116), .A3(new_n816_), .A4(new_n842_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n820_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n355_), .A2(new_n848_), .A3(new_n273_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n355_), .B2(new_n273_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n283_), .A2(new_n273_), .A3(new_n271_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n328_), .A2(new_n347_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n347_), .B1(new_n344_), .B2(new_n328_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n290_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n289_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n847_), .A2(new_n851_), .B1(new_n852_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n839_), .B1(new_n859_), .B2(new_n656_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n846_), .A2(new_n820_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n815_), .B2(KEYINPUT115), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT116), .B1(new_n862_), .B2(new_n842_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n851_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n852_), .A2(new_n858_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n656_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(KEYINPUT57), .A3(new_n867_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n838_), .A2(new_n860_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n281_), .A2(new_n284_), .A3(new_n744_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n281_), .A2(KEYINPUT112), .A3(new_n284_), .A4(new_n744_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n870_), .B1(new_n875_), .B2(new_n696_), .ZN(new_n876_));
  AOI211_X1 g675(.A(KEYINPUT54), .B(new_n645_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n877_));
  OAI22_X1  g676(.A1(new_n869_), .A2(new_n655_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n664_), .A2(new_n524_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n421_), .A2(new_n567_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n806_), .B1(new_n878_), .B2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n645_), .B1(new_n831_), .B2(KEYINPUT58), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n831_), .A2(KEYINPUT117), .A3(KEYINPUT58), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n656_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(KEYINPUT57), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n655_), .B1(new_n890_), .B2(new_n860_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n875_), .A2(new_n696_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT54), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n875_), .A2(new_n870_), .A3(new_n696_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n881_), .A2(KEYINPUT59), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n883_), .A2(new_n898_), .A3(new_n356_), .ZN(new_n899_));
  INV_X1    g698(.A(G113gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n878_), .A2(new_n882_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n355_), .A2(new_n900_), .ZN(new_n902_));
  OAI22_X1  g701(.A1(new_n899_), .A2(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1340gat));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904_));
  INV_X1    g703(.A(G120gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n838_), .A2(new_n860_), .A3(new_n868_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n893_), .A2(new_n894_), .B1(new_n614_), .B2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT59), .B1(new_n907_), .B2(new_n881_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n743_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n868_), .A2(new_n834_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n889_), .A2(KEYINPUT57), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n614_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n909_), .B1(new_n913_), .B2(new_n896_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n905_), .B1(new_n908_), .B2(new_n914_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n905_), .A2(KEYINPUT60), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n905_), .B1(new_n909_), .B2(KEYINPUT60), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n878_), .A2(new_n882_), .A3(new_n916_), .A4(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n904_), .B1(new_n915_), .B2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n743_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G120gat), .B1(new_n883_), .B2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(KEYINPUT119), .A3(new_n918_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n920_), .A2(new_n923_), .ZN(G1341gat));
  OAI21_X1  g723(.A(new_n401_), .B1(new_n901_), .B2(new_n614_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  OAI211_X1 g726(.A(KEYINPUT120), .B(new_n401_), .C1(new_n901_), .C2(new_n614_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n883_), .A2(new_n898_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n614_), .A2(new_n401_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n927_), .A2(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(G1342gat));
  XOR2_X1   g730(.A(KEYINPUT121), .B(G134gat), .Z(new_n932_));
  NOR2_X1   g731(.A1(new_n696_), .A2(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n878_), .A2(new_n656_), .A3(new_n882_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n929_), .A2(new_n933_), .B1(new_n934_), .B2(new_n403_), .ZN(G1343gat));
  NOR2_X1   g734(.A1(new_n593_), .A2(new_n420_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n893_), .A2(new_n894_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n906_), .A2(new_n614_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n664_), .A2(new_n567_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n940_), .A2(new_n355_), .A3(new_n941_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT122), .B(G141gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1344gat));
  NAND3_X1  g743(.A1(new_n940_), .A2(new_n743_), .A3(new_n941_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT123), .B(G148gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1345gat));
  NAND4_X1  g746(.A1(new_n878_), .A2(new_n655_), .A3(new_n936_), .A4(new_n941_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(KEYINPUT124), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n940_), .A2(new_n950_), .A3(new_n655_), .A4(new_n941_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT61), .B(G155gat), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n949_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n949_), .B2(new_n951_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1346gat));
  NAND2_X1  g754(.A1(new_n940_), .A2(new_n941_), .ZN(new_n956_));
  OAI21_X1  g755(.A(G162gat), .B1(new_n956_), .B2(new_n696_), .ZN(new_n957_));
  OR2_X1    g756(.A1(new_n867_), .A2(G162gat), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n956_), .B2(new_n958_), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n596_), .A2(new_n651_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n420_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n524_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n913_), .A2(new_n962_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(KEYINPUT125), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n913_), .A2(new_n965_), .A3(new_n962_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n966_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(KEYINPUT22), .B(G169gat), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n967_), .A2(new_n355_), .A3(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(G169gat), .B1(new_n963_), .B2(new_n356_), .ZN(new_n970_));
  AND2_X1   g769(.A1(new_n970_), .A2(KEYINPUT62), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n970_), .A2(KEYINPUT62), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n969_), .B1(new_n971_), .B2(new_n972_), .ZN(G1348gat));
  NAND2_X1  g772(.A1(new_n967_), .A2(new_n743_), .ZN(new_n974_));
  INV_X1    g773(.A(G176gat), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n907_), .A2(new_n524_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n909_), .A2(new_n975_), .A3(new_n961_), .ZN(new_n977_));
  AOI22_X1  g776(.A1(new_n974_), .A2(new_n975_), .B1(new_n976_), .B2(new_n977_), .ZN(G1349gat));
  INV_X1    g777(.A(G183gat), .ZN(new_n979_));
  NAND4_X1  g778(.A1(new_n976_), .A2(new_n655_), .A3(new_n420_), .A4(new_n960_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n614_), .A2(new_n377_), .ZN(new_n981_));
  AOI22_X1  g780(.A1(new_n979_), .A2(new_n980_), .B1(new_n967_), .B2(new_n981_), .ZN(G1350gat));
  NAND3_X1  g781(.A1(new_n967_), .A2(new_n656_), .A3(new_n378_), .ZN(new_n983_));
  INV_X1    g782(.A(G190gat), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n696_), .B1(new_n964_), .B2(new_n966_), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n983_), .B1(new_n984_), .B2(new_n985_), .ZN(G1351gat));
  NAND3_X1  g785(.A1(new_n878_), .A2(new_n936_), .A3(new_n960_), .ZN(new_n987_));
  INV_X1    g786(.A(new_n987_), .ZN(new_n988_));
  NAND4_X1  g787(.A1(new_n988_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n355_), .ZN(new_n989_));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n990_));
  NAND4_X1  g789(.A1(new_n878_), .A2(new_n355_), .A3(new_n936_), .A4(new_n960_), .ZN(new_n991_));
  INV_X1    g790(.A(G197gat), .ZN(new_n992_));
  OAI21_X1  g791(.A(new_n990_), .B1(new_n991_), .B2(new_n992_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n991_), .A2(new_n992_), .ZN(new_n994_));
  AND3_X1   g793(.A1(new_n989_), .A2(new_n993_), .A3(new_n994_), .ZN(G1352gat));
  NOR2_X1   g794(.A1(new_n987_), .A2(new_n909_), .ZN(new_n996_));
  XOR2_X1   g795(.A(KEYINPUT127), .B(G204gat), .Z(new_n997_));
  XNOR2_X1  g796(.A(new_n996_), .B(new_n997_), .ZN(G1353gat));
  XOR2_X1   g797(.A(KEYINPUT63), .B(G211gat), .Z(new_n999_));
  NAND3_X1  g798(.A1(new_n988_), .A2(new_n655_), .A3(new_n999_), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1001_));
  OAI21_X1  g800(.A(new_n1001_), .B1(new_n987_), .B2(new_n614_), .ZN(new_n1002_));
  AND2_X1   g801(.A1(new_n1000_), .A2(new_n1002_), .ZN(G1354gat));
  OAI21_X1  g802(.A(G218gat), .B1(new_n987_), .B2(new_n696_), .ZN(new_n1004_));
  OR2_X1    g803(.A1(new_n867_), .A2(G218gat), .ZN(new_n1005_));
  OAI21_X1  g804(.A(new_n1004_), .B1(new_n987_), .B2(new_n1005_), .ZN(G1355gat));
endmodule


