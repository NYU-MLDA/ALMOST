//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203_));
  OAI21_X1  g002(.A(G169gat), .B1(new_n203_), .B2(KEYINPUT84), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT84), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT22), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT85), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT85), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n204_), .A2(new_n207_), .A3(new_n212_), .A4(new_n208_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT86), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n210_), .A2(new_n216_), .A3(new_n211_), .A4(new_n213_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT83), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n221_), .B2(new_n218_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT87), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT25), .B(G183gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT26), .B(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n211_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n206_), .A2(new_n208_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT24), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n228_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n220_), .A2(new_n218_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT83), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n220_), .B(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n236_), .B2(new_n218_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n230_), .A2(KEYINPUT24), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n224_), .A2(new_n225_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n225_), .B1(new_n224_), .B2(new_n240_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n202_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n224_), .A2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT87), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n224_), .A2(new_n225_), .A3(new_n240_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT30), .A3(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G99gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G15gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT88), .B(G43gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  NAND4_X1  g052(.A1(new_n243_), .A2(new_n247_), .A3(KEYINPUT89), .A4(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n243_), .A2(new_n247_), .A3(KEYINPUT89), .ZN(new_n255_));
  INV_X1    g054(.A(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT89), .B1(new_n243_), .B2(new_n247_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n254_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT90), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT91), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n258_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT91), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(KEYINPUT90), .A3(new_n264_), .A4(new_n254_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n260_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G113gat), .B(G120gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT31), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n261_), .A2(new_n265_), .A3(new_n267_), .A4(new_n271_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT104), .ZN(new_n276_));
  XOR2_X1   g075(.A(G8gat), .B(G36gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(G92gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT18), .B(G64gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT19), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT20), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n222_), .A2(new_n239_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT101), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n232_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n236_), .A2(KEYINPUT23), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n238_), .B1(new_n288_), .B2(new_n219_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT101), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n237_), .B1(G183gat), .B2(G190gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT22), .B(G169gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n229_), .B1(new_n292_), .B2(new_n208_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n287_), .A2(new_n290_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G197gat), .B(G204gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT21), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G211gat), .B(G218gat), .Z(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n295_), .A2(new_n296_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n284_), .B1(new_n294_), .B2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n241_), .A2(new_n242_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n283_), .B(new_n304_), .C1(new_n305_), .C2(new_n303_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n245_), .A2(new_n303_), .A3(new_n246_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n291_), .A2(new_n293_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n233_), .B1(new_n289_), .B2(KEYINPUT101), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n285_), .A2(new_n286_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n284_), .B1(new_n311_), .B2(new_n302_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n283_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n306_), .B1(new_n313_), .B2(KEYINPUT102), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT102), .ZN(new_n315_));
  AOI211_X1 g114(.A(new_n315_), .B(new_n283_), .C1(new_n307_), .C2(new_n312_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n280_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n241_), .A2(new_n242_), .A3(new_n302_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n312_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n282_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n315_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n313_), .A2(KEYINPUT102), .ZN(new_n322_));
  INV_X1    g121(.A(new_n280_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n306_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT103), .B(KEYINPUT0), .Z(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G57gat), .B(G85gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n270_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT94), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n334_));
  INV_X1    g133(.A(G141gat), .ZN(new_n335_));
  INV_X1    g134(.A(G148gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n336_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(KEYINPUT92), .A2(G141gat), .A3(G148gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(KEYINPUT1), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(KEYINPUT1), .ZN(new_n343_));
  INV_X1    g142(.A(G155gat), .ZN(new_n344_));
  INV_X1    g143(.A(G162gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n342_), .B1(new_n347_), .B2(KEYINPUT93), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT93), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n349_), .A3(new_n346_), .ZN(new_n350_));
  AOI211_X1 g149(.A(new_n333_), .B(new_n340_), .C1(new_n348_), .C2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(G155gat), .B2(G162gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT93), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n342_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n340_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT94), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n351_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n338_), .A2(KEYINPUT3), .ZN(new_n361_));
  OR3_X1    g160(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT2), .B1(new_n339_), .B2(KEYINPUT95), .ZN(new_n363_));
  NAND2_X1  g162(.A1(KEYINPUT95), .A2(KEYINPUT2), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n364_), .A2(KEYINPUT92), .B1(G141gat), .B2(G148gat), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n361_), .B(new_n362_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n346_), .A2(new_n341_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT96), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT96), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(new_n370_), .A3(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n332_), .B1(new_n360_), .B2(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n343_), .A2(new_n349_), .A3(new_n346_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n349_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n342_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n333_), .B1(new_n376_), .B2(new_n340_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n357_), .A2(KEYINPUT94), .A3(new_n358_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n371_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n370_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n382_), .A3(new_n270_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n373_), .A2(KEYINPUT4), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n382_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n332_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n331_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n331_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n373_), .B2(new_n383_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n330_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT33), .B(new_n330_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n373_), .A2(new_n389_), .A3(new_n383_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n330_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n384_), .A2(new_n331_), .A3(new_n387_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n393_), .A2(new_n394_), .A3(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n276_), .B1(new_n325_), .B2(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n393_), .A2(new_n394_), .A3(new_n399_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(KEYINPUT104), .A3(new_n324_), .A4(new_n317_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n323_), .A2(KEYINPUT32), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n321_), .A2(new_n322_), .A3(new_n306_), .A4(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT105), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n384_), .A2(new_n387_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n389_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n390_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n396_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT106), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT106), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n409_), .A2(new_n413_), .A3(new_n396_), .A4(new_n410_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n391_), .A3(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n311_), .B2(new_n302_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n245_), .A2(new_n246_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n302_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n320_), .A2(new_n315_), .B1(new_n418_), .B2(new_n283_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n419_), .A2(KEYINPUT105), .A3(new_n322_), .A4(new_n404_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n307_), .A2(new_n283_), .A3(new_n312_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(new_n418_), .B2(new_n283_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(KEYINPUT32), .A3(new_n323_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n407_), .A2(new_n415_), .A3(new_n420_), .A4(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n401_), .A2(new_n403_), .A3(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n360_), .A2(new_n372_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n302_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G228gat), .ZN(new_n429_));
  INV_X1    g228(.A(G233gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT97), .B1(new_n428_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n303_), .B1(new_n385_), .B2(KEYINPUT29), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT97), .ZN(new_n434_));
  INV_X1    g233(.A(new_n431_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n428_), .A2(KEYINPUT98), .A3(new_n431_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT98), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n432_), .A2(new_n436_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G78gat), .B(G106gat), .Z(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT100), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n441_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n385_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G22gat), .B(G50gat), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n446_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n442_), .A2(new_n443_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n432_), .A2(new_n436_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n437_), .A2(new_n439_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT100), .ZN(new_n457_));
  INV_X1    g256(.A(new_n441_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(KEYINPUT99), .A3(new_n458_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n452_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n456_), .A2(new_n458_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT99), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n443_), .A3(new_n465_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n453_), .A2(new_n459_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n425_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n442_), .A2(new_n459_), .A3(new_n443_), .A4(new_n452_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n466_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(new_n462_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n415_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT27), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n325_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n422_), .B2(new_n280_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n324_), .A2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .A4(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n275_), .B1(new_n468_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n273_), .A2(new_n472_), .A3(new_n274_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n463_), .A2(new_n466_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n480_), .A2(new_n474_), .A3(new_n469_), .A4(new_n476_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G29gat), .B(G36gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(G43gat), .B(G50gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G43gat), .B(G50gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493_));
  INV_X1    g292(.A(G1gat), .ZN(new_n494_));
  INV_X1    g293(.A(G8gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G8gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n497_), .A2(new_n498_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n492_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n492_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n485_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT78), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT78), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n506_), .B(new_n485_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n500_), .A2(new_n499_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n488_), .A2(new_n491_), .A3(KEYINPUT15), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT15), .B1(new_n488_), .B2(new_n491_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(new_n501_), .A3(new_n484_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT79), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT79), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n511_), .A2(new_n501_), .A3(new_n514_), .A4(new_n484_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n505_), .A2(new_n507_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G113gat), .B(G141gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G169gat), .B(G197gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n516_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(KEYINPUT82), .A3(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n516_), .A2(KEYINPUT82), .A3(new_n524_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G204gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT5), .B(G176gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT73), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G71gat), .B(G78gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT71), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n538_), .B2(KEYINPUT11), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n537_), .A2(KEYINPUT71), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n537_), .A2(KEYINPUT71), .ZN(new_n541_));
  OR3_X1    g340(.A1(new_n540_), .A2(new_n541_), .A3(KEYINPUT11), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(KEYINPUT11), .A3(new_n536_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(KEYINPUT69), .A2(G99gat), .A3(G106gat), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT70), .ZN(new_n551_));
  NAND3_X1  g350(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(new_n556_), .A3(new_n549_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G85gat), .B(G92gat), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n559_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n554_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(KEYINPUT68), .A3(new_n552_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT68), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n563_), .B1(new_n569_), .B2(new_n550_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n560_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT10), .B(G99gat), .Z(new_n573_));
  INV_X1    g372(.A(G106gat), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(KEYINPUT64), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT64), .B1(new_n573_), .B2(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n568_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT65), .B(G92gat), .ZN(new_n578_));
  OAI21_X1  g377(.A(G85gat), .B1(new_n578_), .B2(KEYINPUT9), .ZN(new_n579_));
  NAND2_X1  g378(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT66), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT67), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n581_), .A2(KEYINPUT67), .A3(new_n584_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n577_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n545_), .B1(new_n572_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n588_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n577_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n558_), .A2(new_n561_), .B1(new_n570_), .B2(new_n560_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n543_), .A2(new_n544_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT72), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(G230gat), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n430_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n593_), .A2(new_n594_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(KEYINPUT72), .A3(new_n545_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n590_), .A2(new_n596_), .A3(KEYINPUT12), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n606_), .A3(new_n545_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n600_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n535_), .B1(new_n604_), .B2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n605_), .A2(new_n607_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n534_), .B(new_n603_), .C1(new_n610_), .C2(new_n600_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n609_), .A2(new_n611_), .A3(KEYINPUT13), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT13), .B1(new_n609_), .B2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n483_), .A2(new_n529_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n508_), .A2(G231gat), .A3(G233gat), .ZN(new_n617_));
  INV_X1    g416(.A(G231gat), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n500_), .B(new_n499_), .C1(new_n618_), .C2(new_n430_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n545_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(G211gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT16), .B(G183gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n625_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(KEYINPUT76), .A4(KEYINPUT17), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n595_), .A2(new_n619_), .A3(new_n617_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n621_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n626_), .A2(new_n627_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n628_), .B1(new_n633_), .B2(KEYINPUT17), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n621_), .B2(new_n630_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT77), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT77), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n621_), .A2(new_n630_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n637_), .B(new_n631_), .C1(new_n638_), .C2(new_n634_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G190gat), .B(G218gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n641_), .B(new_n642_), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT36), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n601_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n593_), .A2(new_n594_), .A3(new_n492_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n647_));
  NAND2_X1  g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT35), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT75), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n646_), .A3(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n649_), .A2(new_n650_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n652_), .A2(new_n653_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n644_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n652_), .A2(new_n653_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT36), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n643_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n658_), .A2(new_n661_), .A3(new_n654_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT37), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n616_), .A2(new_n640_), .A3(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n494_), .A3(new_n415_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT38), .ZN(new_n667_));
  INV_X1    g466(.A(new_n663_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n631_), .B1(new_n638_), .B2(new_n634_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n616_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n616_), .A2(KEYINPUT107), .A3(new_n670_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n673_), .A2(new_n415_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n667_), .B1(new_n494_), .B2(new_n675_), .ZN(G1324gat));
  NAND2_X1  g475(.A1(new_n474_), .A2(new_n476_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n665_), .A2(new_n495_), .A3(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n616_), .A2(new_n677_), .A3(new_n670_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G8gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G8gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(G1325gat));
  NAND3_X1  g484(.A1(new_n673_), .A2(new_n275_), .A3(new_n674_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G15gat), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT41), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT41), .ZN(new_n689_));
  INV_X1    g488(.A(G15gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n665_), .A2(new_n690_), .A3(new_n275_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n689_), .A3(new_n691_), .ZN(G1326gat));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n665_), .A2(new_n693_), .A3(new_n471_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n673_), .A2(new_n471_), .A3(new_n674_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(new_n696_), .A3(G22gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(G22gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1327gat));
  NOR2_X1   g498(.A1(new_n663_), .A2(new_n640_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n616_), .A2(new_n700_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n701_), .A2(G29gat), .A3(new_n472_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT37), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n663_), .B(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n615_), .A2(new_n529_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n640_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT43), .B(new_n704_), .C1(new_n478_), .C2(new_n482_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .A4(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n640_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n714_), .A2(KEYINPUT44), .A3(new_n708_), .A4(new_n710_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n415_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G29gat), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n716_), .A2(new_n717_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n702_), .B1(new_n719_), .B2(new_n720_), .ZN(G1328gat));
  NAND3_X1  g520(.A1(new_n713_), .A2(new_n677_), .A3(new_n715_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G36gat), .ZN(new_n723_));
  INV_X1    g522(.A(new_n677_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(G36gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n616_), .A2(new_n700_), .A3(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT45), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n723_), .A2(KEYINPUT46), .A3(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1329gat));
  NAND4_X1  g531(.A1(new_n713_), .A2(new_n715_), .A3(G43gat), .A4(new_n275_), .ZN(new_n733_));
  INV_X1    g532(.A(G43gat), .ZN(new_n734_));
  INV_X1    g533(.A(new_n275_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n701_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1330gat));
  NAND3_X1  g538(.A1(new_n713_), .A2(new_n471_), .A3(new_n715_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(G50gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G50gat), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n467_), .A2(G50gat), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT111), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n742_), .A2(new_n743_), .B1(new_n701_), .B2(new_n745_), .ZN(G1331gat));
  INV_X1    g545(.A(new_n529_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n483_), .A2(new_n747_), .A3(new_n614_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n748_), .A2(new_n663_), .A3(new_n640_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(G57gat), .A3(new_n415_), .ZN(new_n750_));
  INV_X1    g549(.A(G57gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n748_), .A2(new_n640_), .A3(new_n664_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n472_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n754_), .B2(new_n753_), .ZN(G1332gat));
  OR3_X1    g555(.A1(new_n752_), .A2(G64gat), .A3(new_n724_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n749_), .A2(new_n677_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(G64gat), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n758_), .B2(G64gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n761_), .B2(new_n762_), .ZN(G1333gat));
  INV_X1    g562(.A(G71gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n749_), .B2(new_n275_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n765_), .A2(new_n766_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n275_), .A2(new_n764_), .ZN(new_n770_));
  OAI22_X1  g569(.A1(new_n768_), .A2(new_n769_), .B1(new_n752_), .B2(new_n770_), .ZN(G1334gat));
  OR3_X1    g570(.A1(new_n752_), .A2(G78gat), .A3(new_n467_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n749_), .A2(new_n471_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(G78gat), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n773_), .B2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n772_), .B1(new_n776_), .B2(new_n777_), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n614_), .A2(new_n747_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n700_), .B(new_n779_), .C1(new_n478_), .C2(new_n482_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT114), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n415_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n714_), .A2(new_n710_), .A3(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n415_), .A2(G85gat), .ZN(new_n784_));
  OAI22_X1  g583(.A1(new_n782_), .A2(G85gat), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(G1336gat));
  AND2_X1   g585(.A1(new_n781_), .A2(new_n677_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n677_), .A2(new_n578_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT115), .ZN(new_n789_));
  OAI22_X1  g588(.A1(new_n787_), .A2(G92gat), .B1(new_n783_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n783_), .B2(new_n735_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n573_), .A3(new_n275_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n781_), .A2(new_n574_), .A3(new_n471_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n714_), .A2(new_n471_), .A3(new_n710_), .A4(new_n779_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n796_), .B(new_n803_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n525_), .A2(KEYINPUT82), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n516_), .A2(new_n524_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n640_), .B1(new_n809_), .B2(new_n527_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n609_), .A2(new_n611_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT13), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n609_), .A2(new_n611_), .A3(KEYINPUT13), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n529_), .A2(KEYINPUT116), .A3(new_n640_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n812_), .A2(new_n815_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n614_), .A2(KEYINPUT117), .A3(new_n812_), .A4(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n806_), .B1(new_n822_), .B2(new_n664_), .ZN(new_n823_));
  AOI211_X1 g622(.A(KEYINPUT54), .B(new_n704_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT118), .B1(new_n608_), .B2(KEYINPUT55), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n608_), .A2(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n610_), .A2(new_n600_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n608_), .A2(KEYINPUT118), .A3(KEYINPUT55), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n533_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT56), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n484_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n511_), .A2(new_n501_), .A3(new_n485_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n522_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n525_), .A2(new_n835_), .ZN(new_n836_));
  OR3_X1    g635(.A1(new_n604_), .A2(new_n608_), .A3(new_n533_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n533_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n832_), .A2(new_n836_), .A3(new_n837_), .A4(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n664_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n841_), .B2(new_n840_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n832_), .A2(new_n747_), .A3(new_n837_), .A4(new_n839_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n813_), .A2(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n847_), .B2(new_n663_), .ZN(new_n848_));
  AOI211_X1 g647(.A(KEYINPUT57), .B(new_n668_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n843_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n825_), .B1(new_n850_), .B2(new_n669_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n275_), .A2(new_n415_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n481_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n747_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n825_), .B1(new_n850_), .B2(new_n709_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n857_), .ZN(new_n859_));
  OAI22_X1  g658(.A1(new_n855_), .A2(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n747_), .A2(G113gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n856_), .B1(new_n861_), .B2(new_n862_), .ZN(G1340gat));
  OAI21_X1  g662(.A(G120gat), .B1(new_n860_), .B2(new_n614_), .ZN(new_n864_));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n614_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n855_), .B(new_n866_), .C1(KEYINPUT60), .C2(new_n865_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n855_), .B2(new_n640_), .ZN(new_n869_));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n669_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n861_), .B2(new_n871_), .ZN(G1342gat));
  AOI21_X1  g671(.A(G134gat), .B1(new_n855_), .B2(new_n668_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n704_), .A2(G134gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n861_), .B2(new_n874_), .ZN(G1343gat));
  NOR2_X1   g674(.A1(new_n275_), .A2(new_n467_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n415_), .A3(new_n724_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n851_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n747_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT119), .B(G141gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n615_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT120), .B(G148gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1345gat));
  NAND2_X1  g683(.A1(new_n878_), .A2(new_n640_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT121), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n878_), .A2(new_n887_), .A3(new_n640_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n886_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1346gat));
  NAND2_X1  g691(.A1(new_n704_), .A2(G162gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT122), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n878_), .A2(new_n894_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n851_), .A2(new_n663_), .A3(new_n877_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(G162gat), .B2(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT123), .ZN(G1347gat));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  INV_X1    g698(.A(new_n479_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n677_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n471_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n858_), .A2(new_n529_), .A3(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n899_), .B1(new_n904_), .B2(new_n206_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n668_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n844_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n640_), .B1(new_n907_), .B2(new_n843_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n747_), .B(new_n902_), .C1(new_n908_), .C2(new_n825_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n904_), .A2(new_n292_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n905_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT124), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n905_), .A2(new_n910_), .A3(new_n914_), .A4(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1348gat));
  NOR2_X1   g715(.A1(new_n858_), .A2(new_n903_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G176gat), .B1(new_n917_), .B2(new_n615_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n851_), .A2(new_n471_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n901_), .A2(new_n208_), .A3(new_n614_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1349gat));
  NAND4_X1  g720(.A1(new_n919_), .A2(new_n677_), .A3(new_n900_), .A4(new_n640_), .ZN(new_n922_));
  INV_X1    g721(.A(G183gat), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n669_), .A2(new_n226_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n922_), .A2(new_n923_), .B1(new_n917_), .B2(new_n924_), .ZN(G1350gat));
  NAND3_X1  g724(.A1(new_n917_), .A2(new_n227_), .A3(new_n668_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n858_), .A2(new_n664_), .A3(new_n903_), .ZN(new_n927_));
  INV_X1    g726(.A(G190gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1351gat));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT125), .B1(new_n876_), .B2(new_n472_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n876_), .A2(KEYINPUT125), .A3(new_n472_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n677_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n851_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n747_), .ZN(new_n936_));
  INV_X1    g735(.A(G197gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n930_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n937_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n935_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n747_), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(G1352gat));
  NAND2_X1  g740(.A1(new_n935_), .A2(new_n615_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g742(.A1(new_n851_), .A2(new_n669_), .A3(new_n934_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  AND2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n944_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n947_), .B1(new_n944_), .B2(new_n945_), .ZN(G1354gat));
  AOI21_X1  g747(.A(G218gat), .B1(new_n935_), .B2(new_n668_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n704_), .A2(G218gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n935_), .B2(new_n950_), .ZN(G1355gat));
endmodule


