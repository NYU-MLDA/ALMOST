//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(KEYINPUT3), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT88), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(KEYINPUT88), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G155gat), .ZN(new_n218_));
  INV_X1    g017(.A(G162gat), .ZN(new_n219_));
  OR3_X1    g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT1), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n218_), .B2(new_n219_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(new_n221_), .C1(G155gat), .C2(G162gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n208_), .A3(new_n206_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n203_), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n225_));
  INV_X1    g024(.A(G22gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n217_), .A2(new_n223_), .A3(KEYINPUT28), .A4(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n226_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n202_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n227_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G197gat), .B(G204gat), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT21), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G197gat), .B(G204gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OR3_X1    g039(.A1(new_n236_), .A2(new_n239_), .A3(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(G228gat), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OR3_X1    g047(.A1(new_n233_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(new_n233_), .B2(new_n243_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n225_), .A2(new_n228_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G22gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(G50gat), .A3(new_n229_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n232_), .A2(new_n255_), .A3(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n249_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n252_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n260_), .A2(new_n261_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(new_n232_), .A3(new_n255_), .A4(new_n258_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268_));
  XOR2_X1   g067(.A(G127gat), .B(G134gat), .Z(new_n269_));
  XOR2_X1   g068(.A(G113gat), .B(G120gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT82), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(G169gat), .A3(G176gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n282_));
  INV_X1    g081(.A(G183gat), .ZN(new_n283_));
  INV_X1    g082(.A(G190gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT23), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(G183gat), .A3(G190gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n282_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(KEYINPUT26), .B(G190gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT80), .B(G183gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT25), .ZN(new_n291_));
  OR2_X1    g090(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n289_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n281_), .B(new_n288_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n287_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(new_n285_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(G190gat), .B2(new_n290_), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT84), .B(G176gat), .Z(new_n302_));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n303_), .A2(new_n304_), .A3(G169gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(G169gat), .B1(new_n303_), .B2(new_n304_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n301_), .A2(new_n278_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G227gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(G71gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G99gat), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n297_), .A2(new_n308_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n297_), .B2(new_n308_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n272_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n308_), .B1(new_n296_), .B2(new_n295_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n312_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n297_), .A2(new_n308_), .A3(new_n312_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n271_), .A3(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G15gat), .B(G43gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT86), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT30), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT31), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n315_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n268_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n324_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n313_), .A2(new_n314_), .A3(new_n272_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n271_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n315_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(KEYINPUT87), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n267_), .A2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT94), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n297_), .A2(new_n243_), .A3(new_n308_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT20), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n282_), .B1(new_n280_), .B2(new_n273_), .ZN(new_n345_));
  XOR2_X1   g144(.A(KEYINPUT25), .B(G183gat), .Z(new_n346_));
  OAI211_X1 g145(.A(new_n300_), .B(new_n345_), .C1(new_n289_), .C2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G169gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n302_), .A2(new_n348_), .B1(new_n277_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n285_), .A2(new_n287_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(G183gat), .B2(G190gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n350_), .B(new_n352_), .C1(new_n349_), .C2(new_n277_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n344_), .B1(new_n354_), .B2(new_n242_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n343_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n316_), .A2(new_n242_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n347_), .A2(new_n353_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n344_), .B1(new_n363_), .B2(new_n243_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n364_), .A3(new_n359_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n342_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n356_), .A2(new_n360_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n359_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n366_), .B1(new_n369_), .B2(new_n342_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G1gat), .B(G29gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT98), .B(G85gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT0), .B(G57gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT97), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n224_), .A2(new_n272_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT96), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n217_), .A2(new_n223_), .A3(new_n271_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n217_), .A2(new_n223_), .A3(new_n271_), .A4(KEYINPUT96), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT4), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n379_), .A2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n378_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n382_), .A2(new_n383_), .B1(G225gat), .B2(G233gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n375_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n375_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT99), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n391_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n370_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(KEYINPUT33), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n384_), .A2(new_n386_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n376_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n382_), .A2(new_n383_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n377_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n375_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(new_n390_), .B2(KEYINPUT33), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n361_), .A2(new_n341_), .A3(new_n365_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n361_), .A2(new_n365_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n341_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n361_), .A2(new_n365_), .A3(KEYINPUT95), .A4(new_n341_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n397_), .A2(new_n403_), .A3(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n335_), .B1(new_n395_), .B2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n327_), .A2(new_n333_), .A3(new_n265_), .A4(new_n263_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n331_), .A2(new_n332_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n266_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n394_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT100), .B1(new_n418_), .B2(new_n392_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT100), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n393_), .A2(new_n420_), .A3(new_n394_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n367_), .A2(new_n368_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n408_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n404_), .A2(KEYINPUT27), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n411_), .A2(new_n422_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n417_), .A2(new_n419_), .A3(new_n421_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n413_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G29gat), .B(G36gat), .Z(new_n430_));
  XOR2_X1   g229(.A(G43gat), .B(G50gat), .Z(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G29gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G43gat), .B(G50gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT15), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n432_), .A2(KEYINPUT15), .A3(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G22gat), .ZN(new_n442_));
  INV_X1    g241(.A(G1gat), .ZN(new_n443_));
  INV_X1    g242(.A(G8gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT14), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G8gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n441_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n436_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n436_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n448_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G113gat), .B(G141gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT79), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G169gat), .B(G197gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n462_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n453_), .A2(new_n457_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT68), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT67), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(G71gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n310_), .A2(KEYINPUT67), .ZN(new_n471_));
  OAI21_X1  g270(.A(G78gat), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G64gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n310_), .A2(KEYINPUT67), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(G71gat), .ZN(new_n476_));
  INV_X1    g275(.A(G78gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n472_), .A2(new_n474_), .A3(KEYINPUT11), .A4(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT11), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n477_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n472_), .A2(KEYINPUT11), .A3(new_n478_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n473_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(G106gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .A4(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT66), .ZN(new_n496_));
  XOR2_X1   g295(.A(G85gat), .B(G92gat), .Z(new_n497_));
  AND3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT8), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n497_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(KEYINPUT66), .A3(new_n500_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n504_));
  INV_X1    g303(.A(G85gat), .ZN(new_n505_));
  OR2_X1    g304(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n512_), .A2(new_n513_), .A3(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n492_), .A2(new_n493_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n503_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n479_), .B(new_n485_), .C1(new_n501_), .C2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n485_), .A2(new_n479_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n502_), .A2(KEYINPUT66), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(KEYINPUT8), .A3(new_n522_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n499_), .A2(new_n500_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G230gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT64), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n468_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  AOI211_X1 g329(.A(KEYINPUT68), .B(new_n530_), .C1(new_n519_), .C2(new_n525_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n519_), .A2(KEYINPUT12), .A3(new_n525_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(new_n524_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n479_), .A4(new_n485_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n528_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT70), .ZN(new_n540_));
  XOR2_X1   g339(.A(G176gat), .B(G204gat), .Z(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n540_), .B(new_n541_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n532_), .A2(new_n538_), .A3(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n544_), .A2(new_n547_), .A3(KEYINPUT71), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT71), .B1(new_n544_), .B2(new_n547_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n532_), .B2(new_n538_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n549_), .B1(new_n553_), .B2(KEYINPUT72), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n537_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n552_), .ZN(new_n557_));
  OAI22_X1  g356(.A1(new_n554_), .A2(new_n557_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(KEYINPUT72), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n556_), .B1(new_n555_), .B2(new_n552_), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n559_), .A2(new_n560_), .A3(new_n549_), .A4(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n485_), .A2(new_n479_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n485_), .B2(new_n479_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n576_), .A2(new_n577_), .A3(KEYINPUT75), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n520_), .A2(new_n573_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n575_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n448_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT75), .B1(new_n576_), .B2(new_n577_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n579_), .A3(new_n575_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(new_n450_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n572_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n582_), .A2(KEYINPUT77), .A3(new_n585_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n570_), .A2(new_n571_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n582_), .A2(KEYINPUT77), .A3(new_n585_), .A4(new_n588_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n586_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT78), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AOI211_X1 g393(.A(KEYINPUT78), .B(new_n586_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n440_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n523_), .A2(new_n524_), .A3(new_n436_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT35), .B(new_n597_), .C1(new_n598_), .C2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n441_), .A2(new_n534_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .A4(new_n599_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n601_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n605_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT74), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n601_), .B2(new_n609_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT37), .B1(new_n610_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n601_), .A2(new_n609_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n612_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n601_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n594_), .A2(new_n595_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR4_X1   g423(.A1(new_n429_), .A2(new_n467_), .A3(new_n565_), .A4(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n421_), .A2(new_n419_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n443_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n618_), .A2(new_n620_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n594_), .A2(new_n595_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n429_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n564_), .A2(new_n466_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT101), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(new_n627_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n629_), .B1(new_n443_), .B2(new_n638_), .ZN(G1324gat));
  INV_X1    g438(.A(new_n426_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G8gat), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT102), .A3(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(G8gat), .A3(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n625_), .A2(new_n444_), .A3(new_n640_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n644_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n644_), .A2(KEYINPUT40), .A3(new_n646_), .A4(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n637_), .B2(new_n334_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n625_), .A2(new_n653_), .A3(new_n334_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n655_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT104), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n656_), .A2(new_n661_), .A3(new_n657_), .A4(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1326gat));
  AOI21_X1  g462(.A(new_n226_), .B1(new_n637_), .B2(new_n267_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT42), .Z(new_n665_));
  NAND3_X1  g464(.A1(new_n625_), .A2(new_n226_), .A3(new_n267_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1327gat));
  NOR2_X1   g466(.A1(new_n632_), .A2(new_n630_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(new_n564_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n428_), .A3(new_n466_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n627_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n428_), .A2(new_n622_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n622_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n413_), .B2(new_n427_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT43), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n633_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n636_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT105), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n679_), .C2(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n627_), .A2(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n672_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  NOR2_X1   g486(.A1(new_n426_), .A2(G36gat), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n670_), .A2(KEYINPUT106), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT106), .B1(new_n670_), .B2(new_n689_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT45), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n426_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n694_));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT46), .B(new_n693_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  XNOR2_X1  g499(.A(KEYINPUT107), .B(G43gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n334_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n670_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT108), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n415_), .A2(G43gat), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n685_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n708_), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n704_), .B(new_n710_), .C1(new_n685_), .C2(new_n706_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n671_), .B2(new_n267_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n266_), .A2(new_n202_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n685_), .B2(new_n714_), .ZN(G1331gat));
  NOR2_X1   g514(.A1(new_n564_), .A2(new_n466_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n634_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n626_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n429_), .A2(new_n466_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n624_), .A2(new_n564_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT110), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(KEYINPUT110), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n720_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(G57gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n627_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n719_), .A2(new_n726_), .ZN(G1332gat));
  OAI21_X1  g526(.A(G64gat), .B1(new_n718_), .B2(new_n426_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n426_), .A2(G64gat), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT112), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n724_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1333gat));
  AOI21_X1  g533(.A(new_n310_), .B1(new_n717_), .B2(new_n334_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT49), .Z(new_n736_));
  NAND3_X1  g535(.A1(new_n724_), .A2(new_n310_), .A3(new_n334_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1334gat));
  AOI21_X1  g537(.A(new_n477_), .B1(new_n717_), .B2(new_n267_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n724_), .A2(new_n477_), .A3(new_n267_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1335gat));
  NAND3_X1  g542(.A1(new_n720_), .A2(new_n565_), .A3(new_n668_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n505_), .A3(new_n627_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n633_), .B1(new_n677_), .B2(KEYINPUT43), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n674_), .B(new_n676_), .C1(new_n413_), .C2(new_n427_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(new_n716_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n627_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n751_), .B2(new_n505_), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n745_), .B2(new_n640_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n426_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n750_), .B2(new_n754_), .ZN(G1337gat));
  NOR2_X1   g554(.A1(new_n512_), .A2(new_n513_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n745_), .A2(new_n756_), .A3(new_n415_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n750_), .A2(new_n334_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n487_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n745_), .A2(new_n488_), .A3(new_n267_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n632_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(new_n267_), .A3(new_n678_), .A4(new_n716_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n749_), .A2(KEYINPUT114), .A3(new_n267_), .A4(new_n716_), .ZN(new_n767_));
  AND4_X1   g566(.A1(new_n762_), .A2(new_n766_), .A3(G106gat), .A4(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n488_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n762_), .B1(new_n769_), .B2(new_n767_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n761_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n761_), .C1(new_n768_), .C2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  NAND3_X1  g574(.A1(new_n564_), .A2(new_n623_), .A3(new_n467_), .ZN(new_n776_));
  OR2_X1    g575(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT116), .Z(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n780_), .A3(new_n777_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n449_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n455_), .A2(new_n452_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n462_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n465_), .A2(new_n787_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT118), .Z(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT119), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n533_), .A2(new_n528_), .A3(new_n536_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT117), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n533_), .A2(new_n794_), .A3(new_n528_), .A4(new_n536_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n537_), .A2(KEYINPUT55), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n798_), .B(new_n528_), .C1(new_n533_), .C2(new_n536_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n796_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n552_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n538_), .A2(new_n798_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n799_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n793_), .A4(new_n795_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  INV_X1    g604(.A(new_n552_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n801_), .A2(new_n466_), .A3(new_n549_), .A4(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n789_), .B(new_n809_), .C1(new_n554_), .C2(new_n557_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n791_), .A2(new_n808_), .A3(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT57), .B1(new_n811_), .B2(new_n630_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n801_), .A2(new_n549_), .A3(new_n807_), .A4(new_n789_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n804_), .A2(new_n806_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n818_), .A2(KEYINPUT56), .B1(new_n555_), .B2(new_n548_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n819_), .A2(new_n815_), .A3(new_n807_), .A4(new_n789_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n676_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n812_), .A2(new_n813_), .A3(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n784_), .B1(new_n822_), .B2(new_n632_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n626_), .A2(new_n640_), .A3(new_n416_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n817_), .A2(new_n820_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n622_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT121), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n821_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n811_), .A2(new_n630_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n829_), .A2(new_n831_), .A3(new_n834_), .A4(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n633_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n784_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n838_), .A2(new_n825_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n466_), .B(new_n826_), .C1(new_n839_), .C2(new_n824_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G113gat), .ZN(new_n841_));
  INV_X1    g640(.A(G113gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n842_), .A3(new_n466_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1340gat));
  OAI211_X1 g643(.A(new_n565_), .B(new_n826_), .C1(new_n839_), .C2(new_n824_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(G120gat), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n564_), .A2(KEYINPUT60), .ZN(new_n847_));
  MUX2_X1   g646(.A(new_n847_), .B(KEYINPUT60), .S(G120gat), .Z(new_n848_));
  NAND2_X1  g647(.A1(new_n839_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(G1341gat));
  OAI211_X1 g649(.A(new_n632_), .B(new_n826_), .C1(new_n839_), .C2(new_n824_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G127gat), .ZN(new_n852_));
  INV_X1    g651(.A(G127gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n839_), .A2(new_n853_), .A3(new_n632_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1342gat));
  OAI211_X1 g654(.A(new_n622_), .B(new_n826_), .C1(new_n839_), .C2(new_n824_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G134gat), .ZN(new_n857_));
  INV_X1    g656(.A(G134gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n839_), .A2(new_n858_), .A3(new_n631_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1343gat));
  NAND2_X1  g659(.A1(new_n782_), .A2(new_n783_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n836_), .B2(new_n633_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n414_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n626_), .A2(new_n640_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n466_), .A3(new_n864_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT122), .B(G141gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1344gat));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n565_), .A3(new_n864_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT123), .B(G148gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1345gat));
  NAND3_X1  g669(.A1(new_n863_), .A2(new_n632_), .A3(new_n864_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  AND2_X1   g672(.A1(new_n863_), .A2(new_n864_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n219_), .A3(new_n631_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n874_), .A2(new_n622_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n219_), .ZN(G1347gat));
  AND2_X1   g676(.A1(new_n466_), .A2(new_n348_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n834_), .A2(new_n828_), .A3(new_n835_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n861_), .B1(new_n879_), .B2(new_n633_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n627_), .A2(new_n426_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n334_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n266_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n880_), .A2(new_n881_), .A3(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n883_), .A2(new_n267_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT125), .B1(new_n823_), .B2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n878_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n823_), .A2(new_n466_), .A3(new_n887_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n890_), .A2(G169gat), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n890_), .B2(G169gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n889_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT126), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n889_), .B(new_n896_), .C1(new_n892_), .C2(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1348gat));
  NAND3_X1  g697(.A1(new_n884_), .A2(G176gat), .A3(new_n565_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n862_), .A2(new_n267_), .A3(new_n899_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n886_), .A2(new_n888_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n565_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n902_), .B2(new_n302_), .ZN(G1349gat));
  AND2_X1   g702(.A1(new_n632_), .A2(new_n346_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n290_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n838_), .A2(new_n266_), .A3(new_n632_), .A4(new_n884_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n901_), .A2(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1350gat));
  INV_X1    g706(.A(new_n289_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n901_), .A2(new_n908_), .A3(new_n631_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n901_), .A2(new_n622_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n284_), .ZN(G1351gat));
  NAND3_X1  g710(.A1(new_n863_), .A2(new_n466_), .A3(new_n882_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g712(.A1(new_n863_), .A2(new_n565_), .A3(new_n882_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g714(.A1(new_n863_), .A2(new_n632_), .A3(new_n882_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  AND2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(new_n916_), .B2(new_n917_), .ZN(G1354gat));
  NOR2_X1   g719(.A1(new_n630_), .A2(G218gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n863_), .A2(new_n882_), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n882_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n862_), .A2(new_n414_), .A3(new_n676_), .A4(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n922_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT127), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n922_), .B(new_n928_), .C1(new_n925_), .C2(new_n924_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1355gat));
endmodule


