//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n913_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n206_), .B1(G155gat), .B2(G162gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(G155gat), .A3(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(G155gat), .B2(G162gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n202_), .B(new_n205_), .C1(new_n207_), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n202_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n218_));
  XOR2_X1   g017(.A(G155gat), .B(G162gat), .Z(new_n219_));
  AND3_X1   g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n218_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n210_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT21), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT89), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT89), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT21), .ZN(new_n228_));
  AND2_X1   g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n226_), .B(new_n228_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(G197gat), .A2(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT21), .A3(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT90), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT90), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n231_), .A2(new_n234_), .A3(new_n238_), .A4(new_n235_), .ZN(new_n239_));
  OR3_X1    g038(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT91), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT91), .B1(new_n234_), .B2(new_n235_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n237_), .A2(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(G228gat), .B(G233gat), .C1(new_n224_), .C2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G78gat), .B(G106gat), .Z(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(new_n239_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n240_), .A2(new_n241_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G228gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT88), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n252_), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(KEYINPUT92), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n243_), .A2(new_n245_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n222_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT28), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G22gat), .B(G50gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n245_), .B1(new_n243_), .B2(new_n255_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n257_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n258_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n263_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n256_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n275_));
  INV_X1    g074(.A(G134gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G127gat), .ZN(new_n277_));
  INV_X1    g076(.A(G127gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G134gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G120gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G113gat), .ZN(new_n282_));
  INV_X1    g081(.A(G113gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G120gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n277_), .A2(new_n279_), .A3(new_n282_), .A4(new_n284_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n275_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n277_), .A2(new_n279_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT82), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT83), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  AND4_X1   g090(.A1(new_n277_), .A2(new_n279_), .A3(new_n282_), .A4(new_n284_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT82), .B1(new_n292_), .B2(new_n289_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT83), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n286_), .A2(new_n275_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n291_), .A2(new_n296_), .A3(KEYINPUT31), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT31), .B1(new_n291_), .B2(new_n296_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT84), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT85), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G43gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT80), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G71gat), .ZN(new_n305_));
  INV_X1    g104(.A(G99gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT22), .B(G169gat), .ZN(new_n310_));
  INV_X1    g109(.A(G176gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT79), .B1(new_n313_), .B2(KEYINPUT23), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(KEYINPUT23), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G183gat), .A3(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n314_), .B1(new_n318_), .B2(KEYINPUT79), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n312_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT25), .B(G183gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G190gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n325_), .A2(KEYINPUT24), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT24), .A3(new_n308_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n324_), .A2(new_n318_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G227gat), .A2(G233gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n330_), .B(KEYINPUT81), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT30), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n329_), .B(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n307_), .A2(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n307_), .A2(new_n333_), .B1(new_n299_), .B2(KEYINPUT84), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n300_), .A2(KEYINPUT85), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n302_), .A2(new_n334_), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n335_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n336_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n301_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n222_), .A2(new_n291_), .A3(new_n296_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT97), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n222_), .A2(new_n291_), .A3(new_n296_), .A4(KEYINPUT97), .ZN(new_n345_));
  OAI221_X1 g144(.A(new_n210_), .B1(new_n289_), .B2(new_n292_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n344_), .A2(KEYINPUT4), .A3(new_n345_), .A4(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n222_), .A2(new_n291_), .A3(new_n296_), .A4(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n344_), .A2(new_n350_), .A3(new_n345_), .A4(new_n346_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n274_), .A2(new_n341_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(KEYINPUT95), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n320_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT94), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n312_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n371_), .A2(new_n372_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n324_), .A2(new_n327_), .A3(new_n326_), .ZN(new_n375_));
  OAI22_X1  g174(.A1(new_n373_), .A2(new_n374_), .B1(new_n375_), .B2(new_n319_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT20), .B1(new_n377_), .B2(new_n242_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n250_), .A2(new_n254_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n329_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT19), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n370_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n246_), .A2(KEYINPUT92), .A3(new_n247_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT92), .B1(new_n246_), .B2(new_n247_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n380_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n248_), .B2(new_n376_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(KEYINPUT95), .A3(new_n383_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n385_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT96), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n377_), .A2(new_n394_), .A3(new_n242_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT96), .B1(new_n248_), .B2(new_n376_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n250_), .A2(new_n254_), .A3(new_n329_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n383_), .A2(new_n389_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n369_), .B1(new_n393_), .B2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT95), .B1(new_n391_), .B2(new_n383_), .ZN(new_n402_));
  AOI211_X1 g201(.A(new_n370_), .B(new_n384_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n369_), .B(new_n400_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n365_), .B1(new_n401_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n369_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n386_), .A2(new_n387_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n248_), .B2(new_n376_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT99), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n408_), .A2(new_n329_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n384_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n391_), .A2(new_n383_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n407_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n404_), .A2(new_n415_), .A3(KEYINPUT27), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT100), .B1(new_n406_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n400_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n407_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT27), .B1(new_n419_), .B2(new_n404_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n404_), .A2(new_n415_), .A3(KEYINPUT27), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT100), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n364_), .B1(new_n417_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n341_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n337_), .A2(new_n340_), .A3(KEYINPUT86), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n361_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n359_), .B(new_n429_), .C1(new_n267_), .C2(new_n272_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n420_), .A2(new_n421_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT98), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT98), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n344_), .A2(new_n435_), .A3(new_n345_), .A4(new_n346_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n351_), .A3(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n349_), .A2(new_n350_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n358_), .B1(new_n347_), .B2(new_n438_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n432_), .A2(new_n359_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n353_), .A2(KEYINPUT33), .A3(new_n354_), .A4(new_n358_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n419_), .A2(new_n440_), .A3(new_n404_), .A4(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(KEYINPUT32), .B(new_n369_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n444_), .B(new_n400_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n443_), .B(new_n445_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n274_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n428_), .B1(new_n431_), .B2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n424_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G232gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT35), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT71), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT73), .ZN(new_n456_));
  XOR2_X1   g255(.A(KEYINPUT10), .B(G99gat), .Z(new_n457_));
  INV_X1    g256(.A(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G85gat), .B(G92gat), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT9), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  INV_X1    g261(.A(G92gat), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT9), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT6), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n459_), .A2(new_n461_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT7), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n306_), .A3(new_n458_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT64), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n473_), .A2(new_n470_), .A3(new_n306_), .A4(new_n458_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n466_), .A2(new_n469_), .A3(new_n472_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n460_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT8), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT8), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n475_), .A2(new_n478_), .A3(new_n460_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n468_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G29gat), .B(G36gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G43gat), .B(G50gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT72), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n452_), .A2(KEYINPUT35), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n477_), .A2(new_n479_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n467_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n483_), .B(KEYINPUT15), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n487_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n456_), .B1(new_n486_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT73), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n454_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n486_), .A2(KEYINPUT73), .A3(new_n455_), .A4(new_n491_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G190gat), .B(G218gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT74), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G134gat), .B(G162gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT36), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n496_), .A2(new_n497_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n501_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(KEYINPUT36), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT37), .B1(new_n503_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n496_), .A2(new_n497_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n505_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n496_), .A2(new_n497_), .A3(new_n502_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G127gat), .B(G155gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT16), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G183gat), .B(G211gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT17), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520_));
  INV_X1    g319(.A(G1gat), .ZN(new_n521_));
  INV_X1    g320(.A(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT75), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n526_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT65), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(KEYINPUT65), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT11), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G71gat), .B(G78gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n530_), .A2(KEYINPUT65), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT11), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n531_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT11), .B(new_n535_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n529_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n529_), .A2(new_n542_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n519_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT76), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n540_), .A2(KEYINPUT67), .A3(new_n541_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT67), .B1(new_n540_), .B2(new_n541_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(new_n529_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n529_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n518_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n545_), .A2(new_n546_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n547_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT77), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT77), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n514_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n526_), .B(new_n483_), .Z(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(G229gat), .A3(G233gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n490_), .A2(new_n526_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n526_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n483_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT78), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G113gat), .B(G141gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(G169gat), .B(G197gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n572_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n480_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n542_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n489_), .A2(new_n580_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n551_), .A2(new_n579_), .B1(new_n581_), .B2(new_n578_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n480_), .A2(new_n542_), .B1(G230gat), .B2(G233gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n480_), .A2(new_n542_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT66), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT66), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n480_), .A2(new_n587_), .A3(new_n542_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n581_), .A3(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(G230gat), .A3(G233gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G120gat), .B(G148gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n584_), .A2(new_n590_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(KEYINPUT13), .A3(new_n599_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n602_), .A2(new_n603_), .A3(KEYINPUT69), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT69), .B1(new_n602_), .B2(new_n603_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR4_X1   g405(.A1(new_n449_), .A2(new_n563_), .A3(new_n577_), .A4(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n362_), .A2(G1gat), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n607_), .A2(KEYINPUT101), .A3(new_n608_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n602_), .A2(new_n603_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n576_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n449_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n510_), .A2(new_n512_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n560_), .A3(new_n559_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n362_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n614_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n612_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(new_n417_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n423_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n607_), .A2(new_n522_), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n617_), .A2(new_n629_), .A3(new_n620_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(G8gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n631_), .B2(G8gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  OAI21_X1  g437(.A(G15gat), .B1(new_n621_), .B2(new_n428_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n640_), .ZN(new_n642_));
  INV_X1    g441(.A(G15gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n428_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n607_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(new_n642_), .A3(new_n645_), .ZN(G1326gat));
  OAI21_X1  g445(.A(G22gat), .B1(new_n621_), .B2(new_n273_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT42), .ZN(new_n648_));
  INV_X1    g447(.A(G22gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n607_), .A2(new_n649_), .A3(new_n274_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(G1327gat));
  NOR2_X1   g450(.A1(new_n503_), .A2(new_n507_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n561_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT104), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n449_), .A2(new_n654_), .A3(new_n616_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G29gat), .B1(new_n655_), .B2(new_n363_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n424_), .A2(new_n448_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n514_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT43), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n657_), .A2(new_n661_), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n615_), .A2(new_n561_), .A3(new_n576_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n666_), .A2(G29gat), .A3(new_n363_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n665_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n656_), .B1(new_n667_), .B2(new_n670_), .ZN(G1328gat));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  INV_X1    g471(.A(G36gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n664_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n628_), .B1(new_n674_), .B2(KEYINPUT44), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n670_), .B2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n655_), .A2(new_n673_), .A3(new_n629_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT45), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n655_), .A2(new_n679_), .A3(new_n673_), .A4(new_n629_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n672_), .B1(new_n676_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n666_), .A2(new_n629_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n674_), .A2(KEYINPUT44), .ZN(new_n684_));
  OAI21_X1  g483(.A(G36gat), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n678_), .A2(new_n680_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(KEYINPUT46), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n682_), .A2(new_n687_), .ZN(G1329gat));
  AOI21_X1  g487(.A(G43gat), .B1(new_n655_), .B2(new_n644_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n341_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(G43gat), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n674_), .B2(KEYINPUT44), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n689_), .B1(new_n670_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n695_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n689_), .B(new_n697_), .C1(new_n670_), .C2(new_n693_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1330gat));
  AOI21_X1  g498(.A(G50gat), .B1(new_n655_), .B2(new_n274_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n666_), .A2(G50gat), .A3(new_n274_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n670_), .ZN(G1331gat));
  NOR3_X1   g501(.A1(new_n604_), .A2(new_n619_), .A3(new_n605_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n657_), .A2(new_n703_), .A3(new_n577_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT109), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n657_), .A2(new_n703_), .A3(new_n706_), .A4(new_n577_), .ZN(new_n707_));
  AND4_X1   g506(.A1(G57gat), .A2(new_n705_), .A3(new_n363_), .A4(new_n707_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n563_), .A2(KEYINPUT106), .A3(new_n615_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT106), .B1(new_n563_), .B2(new_n615_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n657_), .A2(new_n577_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT107), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n712_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n709_), .A4(new_n710_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n713_), .A2(new_n363_), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT108), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n717_), .A2(new_n721_), .A3(new_n718_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n708_), .B1(new_n720_), .B2(new_n722_), .ZN(G1332gat));
  NOR2_X1   g522(.A1(new_n628_), .A2(G64gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n713_), .A2(new_n716_), .A3(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n705_), .A2(new_n629_), .A3(new_n707_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(G64gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G64gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT110), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(new_n725_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1333gat));
  AND2_X1   g533(.A1(new_n713_), .A2(new_n716_), .ZN(new_n735_));
  INV_X1    g534(.A(G71gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n644_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n705_), .A2(new_n644_), .A3(new_n707_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(G71gat), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G71gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1334gat));
  INV_X1    g541(.A(G78gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n735_), .A2(new_n743_), .A3(new_n274_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n705_), .A2(new_n274_), .A3(new_n707_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G78gat), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n745_), .A3(G78gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1335gat));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n615_), .A2(new_n562_), .A3(new_n576_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n661_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT43), .B(new_n514_), .C1(new_n424_), .C2(new_n448_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT112), .B(new_n751_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n363_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G85gat), .ZN(new_n759_));
  INV_X1    g558(.A(new_n606_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n712_), .A2(new_n654_), .A3(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n462_), .A3(new_n363_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n750_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n762_), .ZN(new_n764_));
  AOI211_X1 g563(.A(KEYINPUT113), .B(new_n764_), .C1(new_n758_), .C2(G85gat), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n761_), .A2(new_n463_), .A3(new_n629_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n756_), .A2(new_n629_), .A3(new_n757_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n463_), .ZN(G1337gat));
  NAND2_X1  g568(.A1(new_n690_), .A2(new_n457_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n761_), .A2(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n754_), .A2(new_n428_), .ZN(new_n773_));
  OAI211_X1 g572(.A(KEYINPUT114), .B(new_n772_), .C1(new_n773_), .C2(new_n306_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g574(.A1(new_n761_), .A2(new_n458_), .A3(new_n274_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n274_), .B(new_n751_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n776_), .B(new_n782_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1339gat));
  NOR4_X1   g585(.A1(new_n629_), .A2(new_n274_), .A3(new_n362_), .A4(new_n341_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(G230gat), .A2(G233gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n588_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n587_), .B1(new_n480_), .B2(new_n542_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n582_), .A2(new_n791_), .A3(KEYINPUT117), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT67), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n542_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(new_n489_), .A3(KEYINPUT12), .A4(new_n548_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n578_), .B1(new_n480_), .B2(new_n542_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n795_), .A2(new_n586_), .A3(new_n588_), .A4(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n788_), .B1(new_n792_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT118), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n795_), .A2(new_n796_), .A3(new_n583_), .A4(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(KEYINPUT118), .B2(new_n801_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n801_), .A2(KEYINPUT118), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n582_), .A2(new_n583_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n596_), .B1(new_n800_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT56), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n596_), .C1(new_n800_), .C2(new_n807_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n809_), .A2(new_n576_), .A3(new_n599_), .A4(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n565_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n566_), .A2(new_n568_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n570_), .B1(new_n814_), .B2(KEYINPUT119), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(KEYINPUT119), .B2(new_n814_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n575_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n600_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n812_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT57), .B1(new_n820_), .B2(new_n618_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n822_), .B(new_n652_), .C1(new_n812_), .C2(new_n819_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n809_), .A2(new_n599_), .A3(new_n818_), .A4(new_n811_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n514_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n809_), .A2(new_n599_), .A3(new_n811_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT121), .A3(KEYINPUT58), .A4(new_n818_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n825_), .B2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(new_n829_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n562_), .B1(new_n824_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n615_), .A2(new_n577_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT116), .B1(new_n563_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n602_), .A2(new_n603_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n576_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n562_), .A4(new_n514_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(KEYINPUT54), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT116), .B(new_n842_), .C1(new_n563_), .C2(new_n835_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n787_), .B1(new_n834_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n283_), .A3(new_n576_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT122), .B1(new_n834_), .B2(new_n844_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n845_), .A3(new_n849_), .ZN(new_n850_));
  OAI221_X1 g649(.A(new_n787_), .B1(KEYINPUT122), .B2(KEYINPUT59), .C1(new_n834_), .C2(new_n844_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n577_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n847_), .B1(new_n852_), .B2(new_n283_), .ZN(G1340gat));
  OAI21_X1  g652(.A(new_n281_), .B1(new_n615_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n846_), .B(new_n854_), .C1(KEYINPUT60), .C2(new_n281_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n760_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n281_), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n846_), .A2(new_n278_), .A3(new_n562_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n561_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n278_), .ZN(G1342gat));
  NAND3_X1  g659(.A1(new_n846_), .A2(new_n276_), .A3(new_n652_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n514_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n276_), .ZN(G1343gat));
  INV_X1    g662(.A(new_n823_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n820_), .A2(new_n618_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n822_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n833_), .A2(new_n864_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n561_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n841_), .A2(new_n843_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n628_), .A2(new_n274_), .A3(new_n363_), .A4(new_n428_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n870_), .A2(new_n871_), .A3(new_n576_), .A4(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n576_), .B(new_n873_), .C1(new_n834_), .C2(new_n844_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT123), .B(G141gat), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1344gat));
  AOI21_X1  g679(.A(new_n872_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n606_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n562_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n881_), .B2(new_n658_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n834_), .A2(new_n844_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n652_), .A2(new_n887_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n889_), .A2(new_n872_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT125), .B1(new_n888_), .B2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n881_), .A2(new_n887_), .A3(new_n652_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n889_), .A2(new_n514_), .A3(new_n872_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n893_), .B(new_n894_), .C1(new_n895_), .C2(new_n887_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n896_), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n274_), .A2(new_n363_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n628_), .A2(new_n428_), .A3(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n870_), .A2(new_n576_), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G169gat), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n901_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n905_));
  INV_X1    g704(.A(new_n900_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n889_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(new_n310_), .A3(new_n576_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n904_), .A2(new_n905_), .A3(new_n908_), .ZN(G1348gat));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n311_), .A3(new_n837_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n889_), .A2(new_n760_), .A3(new_n906_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n311_), .B2(new_n911_), .ZN(G1349gat));
  NAND3_X1  g711(.A1(new_n870_), .A2(new_n562_), .A3(new_n900_), .ZN(new_n913_));
  MUX2_X1   g712(.A(new_n322_), .B(G183gat), .S(new_n913_), .Z(G1350gat));
  NAND2_X1  g713(.A1(new_n907_), .A2(new_n658_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(G190gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n907_), .A2(new_n323_), .A3(new_n652_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n628_), .A2(new_n430_), .A3(new_n644_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n870_), .A2(new_n576_), .A3(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g720(.A1(new_n870_), .A2(new_n606_), .A3(new_n919_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n923_), .A2(G204gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(G204gat), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT127), .Z(new_n926_));
  AND3_X1   g725(.A1(new_n922_), .A2(new_n924_), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n870_), .A2(new_n562_), .A3(new_n919_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT63), .B(G211gat), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n930_), .B2(new_n933_), .ZN(G1354gat));
  AND2_X1   g733(.A1(new_n870_), .A2(new_n919_), .ZN(new_n935_));
  INV_X1    g734(.A(G218gat), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n935_), .A2(new_n936_), .A3(new_n652_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n935_), .A2(new_n658_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n936_), .ZN(G1355gat));
endmodule


