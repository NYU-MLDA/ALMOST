//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G85gat), .ZN(new_n204_));
  INV_X1    g003(.A(G92gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n208_), .A2(KEYINPUT64), .A3(new_n207_), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT64), .B1(new_n208_), .B2(new_n207_), .ZN(new_n210_));
  OAI221_X1 g009(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT6), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(new_n213_), .C1(G106gat), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n212_), .B(KEYINPUT6), .Z(new_n217_));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n220_));
  AND2_X1   g019(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(new_n220_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  MUX2_X1   g022(.A(new_n220_), .B(new_n222_), .S(new_n223_), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(KEYINPUT66), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n206_), .A2(new_n208_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n216_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  AOI211_X1 g028(.A(KEYINPUT8), .B(new_n227_), .C1(new_n224_), .C2(new_n213_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n215_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G57gat), .B(G64gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT11), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(KEYINPUT11), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n234_), .A2(new_n235_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n231_), .B(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT12), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT12), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n231_), .A2(new_n241_), .A3(new_n237_), .A4(new_n236_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n203_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(new_n202_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G176gat), .B(G204gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT68), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G120gat), .B(G148gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(KEYINPUT69), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT69), .B1(new_n252_), .B2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT13), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT13), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(new_n255_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G127gat), .B(G155gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT16), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G183gat), .B(G211gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G15gat), .B(G22gat), .ZN(new_n266_));
  INV_X1    g065(.A(G1gat), .ZN(new_n267_));
  INV_X1    g066(.A(G8gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT14), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G8gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n270_), .B(new_n271_), .Z(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT75), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G231gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT76), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n238_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n273_), .B(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n265_), .B1(new_n277_), .B2(KEYINPUT17), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(KEYINPUT17), .B2(new_n265_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT77), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n279_), .B(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n258_), .A2(new_n261_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G232gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT35), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G29gat), .B(G36gat), .Z(new_n290_));
  XOR2_X1   g089(.A(G43gat), .B(G50gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n289_), .B1(new_n231_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n292_), .B(KEYINPUT15), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n231_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n231_), .A2(KEYINPUT71), .A3(new_n297_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n296_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n294_), .A2(new_n295_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n288_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n298_), .B1(new_n287_), .B2(new_n286_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n305_), .A2(new_n294_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G190gat), .B(G218gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT73), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G134gat), .B(G162gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT36), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n307_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n304_), .A2(new_n312_), .A3(new_n311_), .A4(new_n306_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(KEYINPUT74), .A3(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT37), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n283_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT78), .ZN(new_n321_));
  INV_X1    g120(.A(new_n272_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n297_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G229gat), .A2(G233gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n272_), .A2(new_n292_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n272_), .B(new_n292_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(G229gat), .A3(G233gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G113gat), .B(G141gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G169gat), .B(G197gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  AND2_X1   g136(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G169gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT22), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT22), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G169gat), .ZN(new_n350_));
  INV_X1    g149(.A(G176gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G169gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(KEYINPUT80), .A3(new_n351_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n346_), .A2(new_n354_), .A3(new_n355_), .A4(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n343_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n343_), .A2(KEYINPUT23), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n347_), .A2(new_n351_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT24), .A3(new_n355_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n363_), .A2(KEYINPUT24), .ZN(new_n365_));
  INV_X1    g164(.A(G183gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT25), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G183gat), .ZN(new_n369_));
  INV_X1    g168(.A(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT26), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT26), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G190gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .A4(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n358_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n358_), .A2(new_n375_), .A3(KEYINPUT81), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G71gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G99gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n380_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G127gat), .B(G134gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n385_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n384_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G15gat), .B(G43gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT82), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT31), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n397_), .B(new_n401_), .Z(new_n402_));
  XOR2_X1   g201(.A(G211gat), .B(G218gat), .Z(new_n403_));
  INV_X1    g202(.A(KEYINPUT21), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G197gat), .B(G204gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT90), .B1(new_n407_), .B2(KEYINPUT21), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n405_), .A2(new_n409_), .A3(new_n404_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n406_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(KEYINPUT91), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT91), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n405_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n412_), .A2(KEYINPUT21), .A3(new_n403_), .A4(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n362_), .A2(new_n342_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n352_), .A2(new_n355_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n365_), .A2(new_n374_), .A3(new_n364_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n340_), .A2(new_n345_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n411_), .A2(new_n415_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n418_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n417_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT19), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT97), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n417_), .A2(new_n426_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT20), .B1(new_n424_), .B2(new_n425_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n358_), .A2(KEYINPUT81), .A3(new_n375_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT81), .B1(new_n358_), .B2(new_n375_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n425_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT93), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n439_), .B(new_n425_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n434_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n430_), .B(new_n433_), .C1(new_n441_), .C2(new_n432_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT18), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT99), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n442_), .A2(KEYINPUT99), .A3(new_n446_), .ZN(new_n450_));
  OAI211_X1 g249(.A(KEYINPUT20), .B(new_n432_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n439_), .B1(new_n380_), .B2(new_n425_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n440_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n446_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n432_), .B1(new_n417_), .B2(new_n426_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n449_), .A2(KEYINPUT27), .A3(new_n450_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT3), .ZN(new_n461_));
  INV_X1    g260(.A(G141gat), .ZN(new_n462_));
  INV_X1    g261(.A(G148gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT2), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G155gat), .A2(G162gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G155gat), .A2(G162gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n471_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n470_), .A2(new_n476_), .A3(KEYINPUT88), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT1), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT1), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n474_), .A2(new_n485_), .A3(new_n475_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n471_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  OR3_X1    g287(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n489_), .A2(new_n490_), .B1(G141gat), .B2(G148gat), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n488_), .A2(KEYINPUT87), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT87), .B1(new_n488_), .B2(new_n491_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n481_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n416_), .B1(new_n494_), .B2(KEYINPUT29), .ZN(new_n495_));
  AND2_X1   g294(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(G228gat), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n498_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G78gat), .B(G106gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n499_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT92), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n494_), .A2(KEYINPUT29), .ZN(new_n505_));
  XOR2_X1   g304(.A(G22gat), .B(G50gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT28), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n505_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n500_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n495_), .A2(new_n498_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n501_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n504_), .A2(new_n508_), .B1(new_n503_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n513_));
  AND4_X1   g312(.A1(new_n513_), .A2(new_n511_), .A3(new_n503_), .A4(new_n508_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n451_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n446_), .B1(new_n516_), .B2(new_n457_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n459_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT94), .B(new_n446_), .C1(new_n516_), .C2(new_n457_), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n388_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n392_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n493_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n488_), .A2(KEYINPUT87), .A3(new_n491_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n525_), .B1(new_n528_), .B2(new_n481_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT4), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n494_), .A2(KEYINPUT95), .A3(new_n396_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT95), .B1(new_n494_), .B2(new_n396_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT96), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n494_), .B2(new_n396_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n528_), .A2(KEYINPUT96), .A3(new_n525_), .A4(new_n481_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n534_), .B1(new_n542_), .B2(KEYINPUT4), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G1gat), .B(G29gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n204_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT0), .B(G57gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n539_), .B(new_n540_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n548_), .B2(new_n533_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n543_), .A2(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n533_), .B(new_n531_), .C1(new_n548_), .C2(new_n530_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n542_), .A2(new_n532_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n547_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n460_), .A2(new_n515_), .A3(new_n522_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n519_), .A2(new_n520_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n543_), .B2(new_n549_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n547_), .B1(new_n542_), .B2(new_n533_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n532_), .B(new_n531_), .C1(new_n548_), .C2(new_n530_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT33), .A4(new_n547_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n556_), .A2(new_n558_), .A3(new_n561_), .A4(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n456_), .A2(KEYINPUT32), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n516_), .A2(new_n457_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n442_), .B2(new_n564_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n515_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n555_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AOI211_X1 g369(.A(KEYINPUT98), .B(new_n515_), .C1(new_n563_), .C2(new_n567_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n402_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n460_), .A2(new_n522_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n515_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n402_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n554_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n336_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n321_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT101), .ZN(new_n579_));
  INV_X1    g378(.A(new_n554_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n267_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n315_), .A2(new_n316_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n336_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n258_), .A2(new_n261_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .A4(new_n282_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G1gat), .B1(new_n590_), .B2(new_n554_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n581_), .A2(new_n582_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n583_), .A2(new_n591_), .A3(new_n592_), .ZN(G1324gat));
  NAND3_X1  g392(.A1(new_n579_), .A2(new_n268_), .A3(new_n573_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n573_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G8gat), .B1(new_n590_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT39), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g398(.A(G15gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n579_), .A2(new_n600_), .A3(new_n575_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G15gat), .B1(new_n590_), .B2(new_n402_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT41), .Z(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(G1326gat));
  INV_X1    g406(.A(new_n515_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(G22gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT103), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n579_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G22gat), .B1(new_n590_), .B2(new_n608_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT42), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(G1327gat));
  NOR3_X1   g413(.A1(new_n588_), .A2(new_n336_), .A3(new_n282_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT43), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n572_), .A2(new_n576_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n617_), .B2(new_n319_), .ZN(new_n618_));
  AOI211_X1 g417(.A(KEYINPUT43), .B(new_n318_), .C1(new_n572_), .C2(new_n576_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT44), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT44), .B(new_n615_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(G29gat), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n554_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n588_), .A2(new_n282_), .A3(new_n584_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n625_), .B2(new_n628_), .ZN(G1328gat));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n622_), .A2(new_n573_), .A3(new_n623_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G36gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n595_), .A2(G36gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n627_), .A2(new_n577_), .A3(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT46), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n630_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n636_), .B1(new_n631_), .B2(G36gat), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n641_), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643_));
  AND4_X1   g442(.A1(new_n643_), .A2(new_n632_), .A3(KEYINPUT46), .A4(new_n637_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n641_), .B2(KEYINPUT46), .ZN(new_n645_));
  OAI22_X1  g444(.A1(new_n640_), .A2(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n638_), .A2(new_n630_), .A3(new_n639_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT105), .B1(new_n641_), .B2(KEYINPUT46), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n651_), .B(KEYINPUT107), .C1(new_n645_), .C2(new_n644_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n652_), .ZN(G1329gat));
  NAND2_X1  g452(.A1(new_n575_), .A2(G43gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n627_), .A2(new_n577_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n402_), .ZN(new_n656_));
  OAI22_X1  g455(.A1(new_n624_), .A2(new_n654_), .B1(G43gat), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g457(.A1(new_n655_), .A2(G50gat), .A3(new_n608_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n624_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(KEYINPUT108), .A3(new_n515_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G50gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT108), .B1(new_n660_), .B2(new_n515_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT109), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(G1331gat));
  AOI21_X1  g465(.A(new_n587_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(new_n588_), .A3(new_n282_), .A4(new_n318_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n554_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(G57gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n588_), .A2(new_n282_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n587_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(G57gat), .A3(new_n580_), .A4(new_n586_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(KEYINPUT110), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(KEYINPUT110), .B2(new_n673_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT111), .Z(G1332gat));
  NAND2_X1  g475(.A1(new_n672_), .A2(new_n586_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G64gat), .B1(new_n677_), .B2(new_n595_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT48), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n595_), .A2(G64gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n668_), .B2(new_n680_), .ZN(G1333gat));
  OAI21_X1  g480(.A(G71gat), .B1(new_n677_), .B2(new_n402_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n402_), .A2(G71gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n668_), .B2(new_n685_), .ZN(G1334gat));
  OAI21_X1  g485(.A(G78gat), .B1(new_n677_), .B2(new_n608_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT50), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n608_), .A2(G78gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n668_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT113), .Z(G1335gat));
  NOR3_X1   g490(.A1(new_n589_), .A2(new_n282_), .A3(new_n584_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n667_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G85gat), .B1(new_n694_), .B2(new_n580_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n618_), .A2(new_n619_), .ZN(new_n696_));
  NOR4_X1   g495(.A1(new_n696_), .A2(new_n587_), .A3(new_n589_), .A4(new_n282_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n554_), .A2(new_n204_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT114), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n695_), .B1(new_n697_), .B2(new_n699_), .ZN(G1336gat));
  NAND3_X1  g499(.A1(new_n694_), .A2(new_n205_), .A3(new_n573_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n697_), .A2(new_n573_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n205_), .ZN(G1337gat));
  NOR3_X1   g502(.A1(new_n693_), .A2(new_n402_), .A3(new_n214_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n697_), .A2(new_n575_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G99gat), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g506(.A(G106gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n694_), .A2(new_n708_), .A3(new_n515_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n697_), .A2(new_n515_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n711_));
  AND4_X1   g510(.A1(KEYINPUT116), .A2(new_n710_), .A3(G106gat), .A4(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(KEYINPUT116), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n708_), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n710_), .A2(new_n714_), .B1(KEYINPUT116), .B2(new_n711_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n709_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g516(.A(KEYINPUT54), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n320_), .B2(new_n336_), .ZN(new_n719_));
  NOR4_X1   g518(.A1(new_n283_), .A2(new_n319_), .A3(KEYINPUT54), .A4(new_n587_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n240_), .A2(new_n242_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n202_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n240_), .A2(new_n203_), .A3(new_n242_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(KEYINPUT55), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT55), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n726_), .A3(new_n202_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT117), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(KEYINPUT117), .A3(new_n727_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n253_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT118), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(KEYINPUT56), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n252_), .A2(new_n587_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n251_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT118), .B1(new_n737_), .B2(new_n731_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n734_), .B(new_n736_), .C1(KEYINPUT56), .C2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n256_), .A2(new_n257_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n323_), .A2(new_n325_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT119), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT119), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n324_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n332_), .B1(new_n327_), .B2(new_n324_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n335_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n740_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n585_), .B1(new_n739_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT57), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n737_), .B2(new_n731_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n735_), .B1(new_n754_), .B2(new_n733_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n732_), .A2(new_n733_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n753_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n755_), .A2(new_n757_), .B1(new_n740_), .B2(new_n748_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n752_), .B1(new_n758_), .B2(new_n585_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT58), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n737_), .A2(new_n753_), .A3(new_n731_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n747_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n763_), .B2(new_n754_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n754_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n765_), .A2(KEYINPUT58), .A3(new_n761_), .A4(new_n762_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n766_), .A3(new_n319_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n751_), .A2(new_n759_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n282_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n721_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n574_), .A2(new_n580_), .A3(new_n575_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(G113gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n587_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT120), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n775_), .A2(KEYINPUT59), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(KEYINPUT59), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n776_), .B(new_n777_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n767_), .B1(new_n750_), .B2(KEYINPUT57), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n758_), .A2(new_n752_), .A3(new_n585_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n769_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n721_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n771_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n783_), .A2(new_n775_), .A3(KEYINPUT59), .A4(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n336_), .B1(new_n778_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n774_), .B1(new_n786_), .B2(new_n773_), .ZN(G1340gat));
  INV_X1    g586(.A(G120gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n589_), .B2(KEYINPUT60), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n772_), .B(new_n789_), .C1(KEYINPUT60), .C2(new_n788_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n589_), .B1(new_n778_), .B2(new_n785_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n788_), .ZN(G1341gat));
  AOI21_X1  g591(.A(G127gat), .B1(new_n772_), .B2(new_n282_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n778_), .A2(new_n785_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n282_), .A2(G127gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT121), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n793_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT122), .ZN(G1342gat));
  INV_X1    g597(.A(G134gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n772_), .A2(new_n799_), .A3(new_n585_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n318_), .B1(new_n778_), .B2(new_n785_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n799_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT123), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n800_), .B(new_n804_), .C1(new_n801_), .C2(new_n799_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1343gat));
  NOR3_X1   g605(.A1(new_n770_), .A2(new_n608_), .A3(new_n575_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n573_), .A2(new_n554_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n336_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(new_n462_), .ZN(G1344gat));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n589_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(new_n463_), .ZN(G1345gat));
  NAND3_X1  g612(.A1(new_n807_), .A2(new_n282_), .A3(new_n808_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT124), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n807_), .A2(new_n816_), .A3(new_n282_), .A4(new_n808_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT61), .B(G155gat), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n815_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1346gat));
  INV_X1    g620(.A(G162gat), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n809_), .A2(new_n822_), .A3(new_n318_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n809_), .B2(new_n584_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT125), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT125), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n826_), .B(new_n822_), .C1(new_n809_), .C2(new_n584_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n823_), .B1(new_n825_), .B2(new_n827_), .ZN(G1347gat));
  NOR2_X1   g627(.A1(new_n595_), .A2(new_n580_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n608_), .A3(new_n575_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n770_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n347_), .B1(new_n831_), .B2(new_n587_), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT62), .Z(new_n833_));
  NAND2_X1  g632(.A1(new_n587_), .A2(new_n356_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT126), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(G1348gat));
  NAND2_X1  g636(.A1(new_n831_), .A2(new_n588_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G176gat), .ZN(G1349gat));
  NOR3_X1   g638(.A1(new_n770_), .A2(new_n769_), .A3(new_n830_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n366_), .A2(KEYINPUT127), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n840_), .A2(new_n367_), .A3(new_n369_), .A4(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(KEYINPUT127), .A2(G183gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n840_), .B2(new_n843_), .ZN(G1350gat));
  NAND4_X1  g643(.A1(new_n831_), .A2(new_n371_), .A3(new_n373_), .A4(new_n585_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n770_), .A2(new_n318_), .A3(new_n830_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n370_), .ZN(G1351gat));
  NAND2_X1  g646(.A1(new_n807_), .A2(new_n829_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n587_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n588_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g652(.A(KEYINPUT63), .B(G211gat), .C1(new_n849_), .C2(new_n282_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT63), .B(G211gat), .Z(new_n855_));
  AND3_X1   g654(.A1(new_n849_), .A2(new_n282_), .A3(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1354gat));
  OR3_X1    g656(.A1(new_n848_), .A2(G218gat), .A3(new_n584_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G218gat), .B1(new_n848_), .B2(new_n318_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1355gat));
endmodule


