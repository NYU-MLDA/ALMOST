//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(new_n202_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211_));
  INV_X1    g010(.A(G1gat), .ZN(new_n212_));
  INV_X1    g011(.A(G8gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G1gat), .B(G8gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n217_), .A2(new_n208_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n217_), .B(new_n208_), .Z(new_n223_));
  INV_X1    g022(.A(new_n221_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G141gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n222_), .A2(new_n225_), .A3(new_n229_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT7), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G106gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT6), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n238_), .A2(new_n241_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245_));
  XOR2_X1   g044(.A(G85gat), .B(G92gat), .Z(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT8), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(new_n249_), .A3(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT70), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n247_), .A2(new_n250_), .A3(KEYINPUT70), .A4(KEYINPUT8), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G92gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT66), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G92gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT65), .B(G85gat), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT9), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT67), .B1(G85gat), .B2(G92gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(KEYINPUT67), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT68), .B1(new_n261_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT9), .ZN(new_n268_));
  AND2_X1   g067(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT66), .B(G92gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n264_), .A2(new_n265_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n267_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n241_), .A2(new_n242_), .ZN(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT10), .B(G99gat), .Z(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT64), .B(G106gat), .Z(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n254_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G71gat), .B(G78gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G57gat), .B(G64gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n284_), .B1(KEYINPUT11), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(KEYINPUT11), .B2(new_n285_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n284_), .A3(KEYINPUT11), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n234_), .B1(new_n283_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n283_), .A2(new_n290_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n252_), .A2(new_n253_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(KEYINPUT71), .A3(new_n289_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(G230gat), .A2(G233gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n293_), .B2(new_n289_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT12), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n283_), .B2(new_n290_), .ZN(new_n300_));
  AOI211_X1 g099(.A(KEYINPUT12), .B(new_n289_), .C1(new_n254_), .C2(new_n282_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n298_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G176gat), .B(G204gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT73), .ZN(new_n305_));
  XOR2_X1   g104(.A(G120gat), .B(G148gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT75), .B1(new_n303_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n297_), .A2(new_n302_), .A3(new_n309_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n297_), .A2(new_n302_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n316_));
  INV_X1    g115(.A(new_n309_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n310_), .A2(new_n314_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n314_), .B1(new_n310_), .B2(new_n318_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT13), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n318_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n316_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n313_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT13), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n319_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT91), .B1(new_n329_), .B2(G204gat), .ZN(new_n330_));
  INV_X1    g129(.A(G204gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n330_), .B1(G197gat), .B2(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n329_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT21), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n331_), .A2(G197gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT92), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n329_), .B2(G204gat), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n334_), .B(new_n335_), .C1(new_n338_), .C2(KEYINPUT21), .ZN(new_n339_));
  INV_X1    g138(.A(new_n335_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(KEYINPUT21), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(KEYINPUT1), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n343_), .B1(new_n345_), .B2(KEYINPUT1), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT86), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n344_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n347_), .B2(new_n346_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT88), .ZN(new_n355_));
  OAI211_X1 g154(.A(G141gat), .B(G148gat), .C1(new_n355_), .C2(KEYINPUT2), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(KEYINPUT2), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT3), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT89), .ZN(new_n362_));
  INV_X1    g161(.A(new_n343_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(new_n345_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n354_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n342_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT90), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G228gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n368_), .A2(G228gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(G233gat), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n367_), .A2(new_n373_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n375_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT93), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n376_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n377_), .B1(new_n382_), .B2(new_n374_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n375_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT93), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n362_), .A2(new_n364_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n353_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT28), .B1(new_n388_), .B2(KEYINPUT29), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT28), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n365_), .A2(new_n390_), .A3(new_n366_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G22gat), .B(G50gat), .Z(new_n393_));
  OR2_X1    g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n381_), .A2(new_n386_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n383_), .A2(new_n384_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n398_), .A2(KEYINPUT93), .A3(new_n394_), .A4(new_n395_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(G183gat), .ZN(new_n401_));
  INV_X1    g200(.A(G190gat), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT23), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT23), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(KEYINPUT81), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(KEYINPUT81), .B2(new_n405_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT80), .ZN(new_n409_));
  INV_X1    g208(.A(G169gat), .ZN(new_n410_));
  INV_X1    g209(.A(G176gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT24), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT24), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT25), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(G183gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT26), .B(G190gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT25), .B(G183gat), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n418_), .B(new_n419_), .C1(new_n420_), .C2(new_n416_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n407_), .A2(new_n413_), .A3(new_n415_), .A4(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT82), .B(G176gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT22), .B(G169gat), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n423_), .A2(new_n424_), .B1(G169gat), .B2(G176gat), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n403_), .B1(KEYINPUT23), .B2(new_n404_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(G183gat), .A2(G190gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n422_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT30), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n429_), .B(KEYINPUT83), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT30), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G43gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G227gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(G15gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n439_), .B(new_n442_), .Z(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n436_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n433_), .A2(new_n435_), .A3(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(KEYINPUT85), .A3(new_n446_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G127gat), .B(G134gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT84), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G120gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT31), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n449_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n455_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n447_), .A2(new_n448_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n400_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT98), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT4), .ZN(new_n462_));
  INV_X1    g261(.A(new_n454_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n388_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n365_), .A2(KEYINPUT95), .A3(new_n463_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT95), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n388_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n454_), .B1(new_n365_), .B2(KEYINPUT95), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n468_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n467_), .B1(new_n472_), .B2(new_n462_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G1gat), .B(G29gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT97), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n472_), .A2(new_n480_), .A3(new_n466_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n470_), .A2(new_n471_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n468_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT97), .B1(new_n484_), .B2(new_n465_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n473_), .B(new_n479_), .C1(new_n481_), .C2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n461_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n480_), .B1(new_n472_), .B2(new_n466_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(KEYINPUT97), .A3(new_n465_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n484_), .A2(KEYINPUT4), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n489_), .A2(new_n490_), .B1(new_n491_), .B2(new_n467_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(KEYINPUT98), .A3(KEYINPUT33), .A4(new_n479_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n342_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n434_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n407_), .B1(G183gat), .B2(G190gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n425_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n426_), .B1(new_n414_), .B2(new_n408_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n420_), .A2(new_n419_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n413_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n497_), .B1(new_n503_), .B2(new_n342_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G226gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT19), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n503_), .A2(new_n342_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT94), .B1(new_n503_), .B2(new_n342_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n431_), .A2(new_n342_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n507_), .A2(new_n497_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n508_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G8gat), .B(G36gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT18), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G64gat), .B(G92gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n508_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n464_), .A2(new_n465_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n484_), .B2(KEYINPUT4), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n478_), .B1(new_n472_), .B2(new_n465_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n523_), .B(new_n524_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n528_), .B1(new_n486_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n494_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n486_), .A2(KEYINPUT101), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT101), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n492_), .A2(new_n534_), .A3(new_n479_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n473_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n478_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n521_), .A2(KEYINPUT32), .ZN(new_n539_));
  INV_X1    g338(.A(new_n507_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n496_), .A2(new_n540_), .A3(new_n504_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n509_), .A2(new_n497_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n540_), .B1(new_n514_), .B2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n539_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT100), .ZN(new_n545_));
  OAI22_X1  g344(.A1(new_n544_), .A2(new_n545_), .B1(new_n517_), .B2(new_n539_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n545_), .B2(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n538_), .A2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n460_), .B1(new_n532_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT27), .B1(new_n523_), .B2(new_n524_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n522_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n552_), .A2(new_n524_), .A3(KEYINPUT27), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n554_), .A2(new_n533_), .A3(new_n535_), .A4(new_n537_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n459_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n400_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n459_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI211_X1 g359(.A(new_n233_), .B(new_n328_), .C1(new_n550_), .C2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT36), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n283_), .A2(new_n210_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT35), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(KEYINPUT76), .A3(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n283_), .A2(new_n208_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n571_), .B2(new_n570_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n570_), .A2(new_n571_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n566_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n581_), .A3(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT77), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT37), .B1(new_n579_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n583_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT16), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT78), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n217_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n289_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n593_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n586_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n561_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n212_), .A3(new_n538_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n602_), .A2(new_n603_), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n583_), .B1(new_n549_), .B2(new_n559_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n599_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n233_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n322_), .A2(new_n610_), .A3(new_n611_), .A4(new_n327_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT103), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT103), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n609_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n212_), .B1(new_n615_), .B2(new_n538_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT104), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n606_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n608_), .A2(new_n617_), .A3(new_n618_), .ZN(G1324gat));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n614_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n550_), .A2(new_n560_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n583_), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT105), .B1(new_n622_), .B2(new_n554_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT105), .ZN(new_n624_));
  INV_X1    g423(.A(new_n554_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n615_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n626_), .A3(G8gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT39), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n623_), .A2(new_n626_), .A3(new_n629_), .A4(G8gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n601_), .A2(new_n213_), .A3(new_n625_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(KEYINPUT40), .A3(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1325gat));
  OAI21_X1  g436(.A(G15gat), .B1(new_n622_), .B2(new_n459_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT41), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(KEYINPUT41), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n601_), .A2(new_n441_), .A3(new_n556_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .ZN(G1326gat));
  OAI21_X1  g441(.A(G22gat), .B1(new_n622_), .B2(new_n400_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT42), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n400_), .A2(G22gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT106), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n601_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(G1327gat));
  NOR2_X1   g447(.A1(new_n583_), .A2(new_n610_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n561_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n538_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n328_), .A2(new_n610_), .A3(new_n233_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n586_), .B1(new_n549_), .B2(new_n559_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n586_), .C1(new_n549_), .C2(new_n559_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT107), .B1(new_n654_), .B2(KEYINPUT43), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n653_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n662_), .A2(G29gat), .A3(new_n538_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n653_), .B(KEYINPUT44), .C1(new_n658_), .C2(new_n659_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n652_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n561_), .A2(new_n666_), .A3(new_n625_), .A4(new_n649_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT45), .Z(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n554_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(new_n664_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n669_), .B(KEYINPUT46), .C1(new_n671_), .C2(new_n666_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n666_), .B1(new_n670_), .B2(new_n664_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n668_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(G1329gat));
  NAND4_X1  g475(.A1(new_n662_), .A2(G43gat), .A3(new_n556_), .A4(new_n664_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n438_), .B1(new_n650_), .B2(new_n459_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1330gat));
  INV_X1    g481(.A(new_n400_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G50gat), .B1(new_n651_), .B2(new_n683_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n662_), .A2(G50gat), .A3(new_n683_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n664_), .ZN(G1331gat));
  NAND2_X1  g485(.A1(new_n328_), .A2(new_n233_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n550_), .B2(new_n560_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n600_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n538_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n610_), .A2(new_n233_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n621_), .A2(new_n328_), .A3(new_n583_), .A4(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n538_), .A2(KEYINPUT109), .A3(G57gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(KEYINPUT109), .B2(G57gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n691_), .B1(new_n695_), .B2(new_n697_), .ZN(G1332gat));
  OAI21_X1  g497(.A(G64gat), .B1(new_n694_), .B2(new_n554_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n554_), .A2(G64gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n689_), .B2(new_n702_), .ZN(G1333gat));
  OAI21_X1  g502(.A(G71gat), .B1(new_n694_), .B2(new_n459_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT49), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n459_), .A2(G71gat), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT111), .Z(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n689_), .B2(new_n707_), .ZN(G1334gat));
  OAI21_X1  g507(.A(G78gat), .B1(new_n694_), .B2(new_n400_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT50), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n400_), .A2(G78gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT112), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n689_), .B2(new_n712_), .ZN(G1335gat));
  NOR2_X1   g512(.A1(new_n687_), .A2(new_n610_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n538_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n271_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n688_), .A2(new_n649_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n538_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1336gat));
  OR3_X1    g521(.A1(new_n715_), .A2(new_n272_), .A3(new_n554_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n255_), .B1(new_n719_), .B2(new_n554_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1337gat));
  OAI21_X1  g524(.A(G99gat), .B1(new_n715_), .B2(new_n459_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n279_), .A3(new_n556_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(G1338gat));
  XNOR2_X1  g529(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n683_), .B(new_n714_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G106gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT52), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n735_), .A3(G106gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n720_), .A2(new_n280_), .A3(new_n683_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n731_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n732_), .A2(new_n735_), .A3(G106gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n735_), .B1(new_n732_), .B2(G106gat), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n738_), .B(new_n731_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n739_), .A2(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(KEYINPUT122), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n611_), .A2(G113gat), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT59), .ZN(new_n747_));
  OAI211_X1 g546(.A(KEYINPUT55), .B(new_n298_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT116), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT12), .B1(new_n293_), .B2(new_n289_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n283_), .A2(new_n299_), .A3(new_n290_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(KEYINPUT55), .A4(new_n298_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n749_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n291_), .B(new_n294_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n756_), .A2(new_n296_), .B1(new_n302_), .B2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n309_), .B1(new_n755_), .B2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(KEYINPUT56), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT56), .ZN(new_n761_));
  AOI211_X1 g560(.A(new_n761_), .B(new_n309_), .C1(new_n755_), .C2(new_n758_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n760_), .A2(new_n762_), .A3(KEYINPUT117), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n755_), .A2(new_n758_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n317_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT117), .A3(new_n761_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n311_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n233_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT118), .B1(new_n763_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n765_), .A2(new_n761_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT117), .B1(new_n759_), .B2(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n766_), .A4(new_n768_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n220_), .A2(KEYINPUT119), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n220_), .A2(KEYINPUT119), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n221_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n229_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n231_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT120), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n325_), .A3(new_n319_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n770_), .A2(new_n775_), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT57), .A3(new_n583_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n760_), .A2(new_n762_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n780_), .A2(KEYINPUT120), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n780_), .A2(KEYINPUT120), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n767_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(KEYINPUT58), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n586_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT58), .B1(new_n785_), .B2(new_n788_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n784_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT57), .B1(new_n783_), .B2(new_n583_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n599_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n586_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n796_), .A2(new_n327_), .A3(new_n322_), .A4(new_n693_), .ZN(new_n797_));
  XOR2_X1   g596(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n795_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n716_), .A2(new_n625_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n557_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n747_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n790_), .A2(new_n791_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n583_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n782_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n773_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(KEYINPUT118), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n808_), .B1(new_n811_), .B2(new_n775_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n807_), .B1(new_n812_), .B2(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(new_n794_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n610_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n747_), .B(new_n805_), .C1(new_n815_), .C2(new_n799_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n804_), .B1(new_n795_), .B2(new_n800_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT121), .A3(new_n747_), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n746_), .B(new_n806_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G113gat), .B1(new_n819_), .B2(new_n611_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n745_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n806_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n746_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n822_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT122), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n828_), .ZN(G1340gat));
  INV_X1    g628(.A(G120gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n818_), .A2(new_n820_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n328_), .B1(new_n819_), .B2(new_n747_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n830_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n328_), .A2(new_n835_), .A3(new_n830_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n835_), .B2(new_n830_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n819_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT123), .B1(new_n834_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n832_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(new_n838_), .C1(new_n842_), .C2(new_n830_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n819_), .B2(new_n610_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n610_), .A2(new_n846_), .A3(G127gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n846_), .B2(G127gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n845_), .B1(new_n824_), .B2(new_n848_), .ZN(G1342gat));
  AOI21_X1  g648(.A(G134gat), .B1(new_n819_), .B2(new_n808_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(KEYINPUT125), .Z(new_n851_));
  AND2_X1   g650(.A1(new_n586_), .A2(G134gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n824_), .B2(new_n852_), .ZN(G1343gat));
  AOI21_X1  g652(.A(new_n558_), .B1(new_n795_), .B2(new_n800_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n802_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n233_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT126), .B(G141gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1344gat));
  INV_X1    g657(.A(new_n328_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n855_), .A2(new_n859_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g660(.A1(new_n855_), .A2(new_n599_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT61), .B(G155gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  OAI21_X1  g663(.A(G162gat), .B1(new_n855_), .B2(new_n796_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n583_), .A2(G162gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n855_), .B2(new_n866_), .ZN(G1347gat));
  NOR3_X1   g666(.A1(new_n557_), .A2(new_n538_), .A3(new_n554_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n801_), .A2(new_n611_), .A3(new_n424_), .A4(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n801_), .A2(new_n611_), .A3(new_n868_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(G169gat), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n872_), .A2(KEYINPUT127), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n870_), .A3(G169gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n872_), .B2(KEYINPUT127), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n869_), .B1(new_n873_), .B2(new_n875_), .ZN(G1348gat));
  NAND2_X1  g675(.A1(new_n801_), .A2(new_n868_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n859_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n411_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n423_), .B2(new_n878_), .ZN(G1349gat));
  NOR2_X1   g679(.A1(new_n877_), .A2(new_n599_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n420_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n401_), .B2(new_n881_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n877_), .B2(new_n796_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n808_), .A2(new_n419_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n877_), .B2(new_n885_), .ZN(G1351gat));
  NAND3_X1  g685(.A1(new_n854_), .A2(new_n716_), .A3(new_n625_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n233_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n329_), .ZN(G1352gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n859_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n331_), .ZN(G1353gat));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n599_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  AND2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n892_), .B2(new_n893_), .ZN(G1354gat));
  OAI21_X1  g695(.A(G218gat), .B1(new_n887_), .B2(new_n796_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n583_), .A2(G218gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n887_), .B2(new_n898_), .ZN(G1355gat));
endmodule


