//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n975_;
  XNOR2_X1  g000(.A(KEYINPUT10), .B(G99gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT64), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT64), .ZN(new_n204_));
  AOI21_X1  g003(.A(G106gat), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT65), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n211_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n207_), .A2(new_n209_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n216_), .A2(G85gat), .A3(G92gat), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(KEYINPUT9), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n205_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  OR3_X1    g024(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n225_), .B1(new_n229_), .B2(KEYINPUT66), .ZN(new_n230_));
  INV_X1    g029(.A(new_n227_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n213_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n213_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n230_), .A2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n231_), .B2(new_n232_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n226_), .A2(new_n241_), .A3(new_n227_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n240_), .B(new_n242_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n223_), .B1(new_n243_), .B2(new_n218_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n222_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G29gat), .B(G36gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G43gat), .B(G50gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT15), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G232gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT34), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(KEYINPUT73), .A3(KEYINPUT35), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n252_), .A2(KEYINPUT35), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n229_), .A2(KEYINPUT66), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n224_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n243_), .A2(new_n218_), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n257_), .A2(new_n258_), .B1(new_n259_), .B2(KEYINPUT8), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n260_), .B2(new_n221_), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT68), .B(new_n222_), .C1(new_n239_), .C2(new_n244_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n248_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT70), .A4(new_n248_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n255_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n252_), .A2(KEYINPUT35), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  AOI211_X1 g071(.A(new_n272_), .B(new_n255_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G190gat), .B(G218gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT36), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT36), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT71), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT72), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(KEYINPUT37), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n274_), .A2(KEYINPUT74), .A3(new_n278_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT74), .B1(new_n274_), .B2(new_n278_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n284_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT37), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G57gat), .B(G64gat), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT11), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(KEYINPUT11), .ZN(new_n294_));
  XOR2_X1   g093(.A(G71gat), .B(G78gat), .Z(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G15gat), .B(G22gat), .ZN(new_n299_));
  INV_X1    g098(.A(G1gat), .ZN(new_n300_));
  INV_X1    g099(.A(G8gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT14), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n298_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT17), .ZN(new_n309_));
  XOR2_X1   g108(.A(G127gat), .B(G155gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G183gat), .B(G211gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n308_), .A2(new_n309_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(KEYINPUT17), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n308_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n291_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n261_), .A2(new_n298_), .A3(new_n262_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n298_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n245_), .A2(KEYINPUT12), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n298_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n322_), .B(new_n324_), .C1(new_n325_), .C2(KEYINPUT12), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G230gat), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n321_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n261_), .A2(new_n262_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n323_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT12), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n322_), .A2(new_n324_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(KEYINPUT69), .A4(new_n327_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n322_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n328_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G120gat), .B(G148gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT5), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G176gat), .B(G204gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n336_), .A2(new_n338_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT13), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(KEYINPUT13), .A3(new_n346_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n320_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G22gat), .B(G50gat), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT83), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(G141gat), .A3(G148gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT2), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT85), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n355_), .A2(new_n359_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(G141gat), .B2(G148gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT3), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT85), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n356_), .A2(new_n358_), .A3(new_n368_), .A4(new_n359_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n361_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n375_), .A3(new_n372_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n356_), .A2(new_n358_), .A3(new_n378_), .A4(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT84), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n356_), .A2(new_n358_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n378_), .A2(new_n379_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT84), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .A4(new_n376_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n374_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT28), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n370_), .A2(new_n373_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n387_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n354_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n353_), .A3(new_n394_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G197gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(G204gat), .ZN(new_n403_));
  INV_X1    g202(.A(G204gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(G197gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT21), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G211gat), .B(G218gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT88), .B1(new_n402_), .B2(G204gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(new_n404_), .A3(G197gat), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n408_), .B(new_n410_), .C1(G197gat), .C2(new_n404_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n406_), .B(new_n407_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n407_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(KEYINPUT21), .A3(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G228gat), .ZN(new_n417_));
  INV_X1    g216(.A(G233gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n387_), .B1(new_n374_), .B2(new_n386_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n390_), .A2(KEYINPUT87), .A3(new_n387_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT90), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n422_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT87), .B1(new_n390_), .B2(new_n387_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .A4(new_n420_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n419_), .B1(new_n421_), .B2(new_n416_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n430_), .A2(new_n435_), .A3(new_n431_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n401_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT91), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n430_), .A2(KEYINPUT91), .A3(new_n435_), .A4(new_n431_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n439_), .A2(new_n401_), .A3(new_n434_), .A4(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n400_), .B1(new_n433_), .B2(new_n432_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n444_), .A2(KEYINPUT92), .A3(new_n440_), .A4(new_n439_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n437_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n374_), .A2(new_n386_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G127gat), .B(G134gat), .Z(new_n448_));
  XOR2_X1   g247(.A(G113gat), .B(G120gat), .Z(new_n449_));
  XOR2_X1   g248(.A(new_n448_), .B(new_n449_), .Z(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n390_), .A2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n451_), .A2(new_n453_), .A3(KEYINPUT4), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n451_), .B2(KEYINPUT4), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT98), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n451_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT99), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n451_), .A2(new_n453_), .A3(KEYINPUT99), .A4(new_n455_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n451_), .A2(new_n453_), .A3(KEYINPUT4), .ZN(new_n464_));
  OR3_X1    g263(.A1(new_n390_), .A2(new_n452_), .A3(KEYINPUT4), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT98), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .A4(new_n456_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G29gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(G85gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT0), .B(G57gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n470_), .B(new_n471_), .Z(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n458_), .A2(new_n463_), .A3(new_n472_), .A4(new_n467_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(KEYINPUT102), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT102), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n468_), .A2(new_n477_), .A3(new_n473_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G169gat), .A2(G176gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT22), .B(G169gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT80), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT22), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT80), .B1(new_n485_), .B2(G169gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(G176gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n481_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(G183gat), .A2(G190gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G183gat), .A2(G190gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n490_), .B1(new_n491_), .B2(KEYINPUT23), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT23), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n493_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(KEYINPUT79), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT79), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G183gat), .A3(G190gat), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(KEYINPUT23), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n488_), .B1(new_n489_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G169gat), .ZN(new_n502_));
  INV_X1    g301(.A(G176gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(KEYINPUT78), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT78), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(G169gat), .B2(G176gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT24), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n504_), .A2(new_n506_), .A3(KEYINPUT24), .A4(new_n480_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT25), .B(G183gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT26), .B(G190gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n493_), .B1(G183gat), .B2(G190gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n496_), .A2(new_n498_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n493_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n501_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G71gat), .B(G99gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(G43gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n519_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G227gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(G15gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT30), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n522_), .A2(new_n526_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT82), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(KEYINPUT82), .A3(new_n528_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n450_), .B(KEYINPUT31), .Z(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n479_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G8gat), .B(G36gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT18), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G64gat), .B(G92gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G226gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT19), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n416_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT20), .B1(new_n519_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n549_), .B1(new_n517_), .B2(new_n489_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT23), .B1(new_n496_), .B2(new_n498_), .ZN(new_n551_));
  OAI221_X1 g350(.A(KEYINPUT95), .B1(G183gat), .B2(G190gat), .C1(new_n551_), .C2(new_n515_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n483_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n482_), .A2(KEYINPUT94), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(new_n503_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n550_), .A2(new_n552_), .A3(new_n556_), .A4(new_n480_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT96), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n482_), .B(new_n553_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n481_), .B1(new_n559_), .B2(new_n503_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n552_), .A4(new_n550_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n514_), .B2(new_n500_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n507_), .A2(new_n508_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n494_), .B(new_n492_), .C1(new_n516_), .C2(new_n493_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(KEYINPUT93), .A4(new_n510_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n558_), .A2(new_n562_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n547_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n548_), .B1(new_n570_), .B2(KEYINPUT97), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n557_), .A2(KEYINPUT96), .B1(new_n564_), .B2(new_n567_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n416_), .B1(new_n572_), .B2(new_n562_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT97), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n546_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n577_));
  AOI211_X1 g376(.A(new_n577_), .B(new_n545_), .C1(new_n519_), .C2(new_n547_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n572_), .A2(new_n416_), .A3(new_n562_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n543_), .B1(new_n576_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n548_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n584_));
  AOI211_X1 g383(.A(KEYINPUT97), .B(new_n416_), .C1(new_n572_), .C2(new_n562_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n545_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n542_), .A3(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT27), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n570_), .A2(KEYINPUT97), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n575_), .A3(new_n583_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n581_), .B1(new_n591_), .B2(new_n545_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n589_), .B1(new_n592_), .B2(new_n542_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n519_), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT20), .B1(new_n594_), .B2(new_n416_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n565_), .A2(new_n566_), .A3(new_n510_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n557_), .A2(new_n416_), .A3(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n545_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n591_), .B2(new_n545_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n543_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n588_), .A2(new_n589_), .B1(new_n593_), .B2(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n446_), .A2(new_n538_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n537_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n443_), .A2(new_n445_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n437_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n576_), .A2(new_n543_), .A3(new_n581_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n542_), .B1(new_n586_), .B2(new_n580_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n589_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n587_), .A3(KEYINPUT27), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n476_), .A2(new_n478_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n603_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n458_), .A2(new_n467_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n472_), .A4(new_n463_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n475_), .A2(KEYINPUT100), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT101), .ZN(new_n620_));
  INV_X1    g419(.A(new_n588_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n616_), .A2(new_n622_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n475_), .A2(new_n617_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n464_), .A2(new_n465_), .A3(new_n455_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n451_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n473_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n624_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n620_), .A2(new_n621_), .A3(new_n623_), .A4(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n599_), .A2(KEYINPUT32), .A3(new_n542_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT32), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n592_), .B1(new_n631_), .B2(new_n543_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n479_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n446_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n602_), .B1(new_n613_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n249_), .A2(new_n305_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n248_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n305_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G229gat), .A2(G233gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT76), .Z(new_n641_));
  XNOR2_X1  g440(.A(new_n305_), .B(new_n637_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n640_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n639_), .A2(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(G113gat), .B(G141gat), .Z(new_n645_));
  XNOR2_X1  g444(.A(G169gat), .B(G197gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT77), .Z(new_n649_));
  OR2_X1    g448(.A1(new_n644_), .A2(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n635_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n352_), .A2(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT103), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(KEYINPUT103), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n655_), .A2(new_n300_), .A3(new_n479_), .A4(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n349_), .A2(new_n350_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n651_), .A3(new_n319_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n288_), .A2(new_n284_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT74), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(new_n279_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n635_), .B2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n446_), .A2(new_n538_), .A3(new_n601_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n629_), .A2(new_n446_), .A3(new_n633_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n537_), .B1(new_n669_), .B2(new_n446_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(KEYINPUT104), .A3(new_n289_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n661_), .B1(new_n666_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G1gat), .B1(new_n674_), .B2(new_n611_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n657_), .A2(new_n658_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n659_), .A2(new_n675_), .A3(new_n676_), .ZN(G1324gat));
  INV_X1    g476(.A(new_n601_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n655_), .A2(new_n301_), .A3(new_n678_), .A4(new_n656_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n673_), .A2(new_n678_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(G8gat), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT39), .B(new_n301_), .C1(new_n673_), .C2(new_n678_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g484(.A1(new_n673_), .A2(new_n603_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G15gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT105), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n686_), .A2(new_n689_), .A3(G15gat), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n688_), .A2(KEYINPUT41), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT41), .B1(new_n688_), .B2(new_n690_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n654_), .A2(G15gat), .A3(new_n537_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(G1326gat));
  OAI21_X1  g493(.A(G22gat), .B1(new_n674_), .B2(new_n446_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT42), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n446_), .A2(G22gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n654_), .B2(new_n697_), .ZN(G1327gat));
  NOR3_X1   g497(.A1(new_n351_), .A2(new_n652_), .A3(new_n319_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n635_), .A2(KEYINPUT43), .A3(new_n291_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n285_), .B1(new_n665_), .B2(KEYINPUT37), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n671_), .B2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n700_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n635_), .B2(new_n291_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n671_), .A2(new_n702_), .A3(new_n701_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(KEYINPUT44), .A3(new_n699_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n707_), .A2(new_n712_), .A3(new_n611_), .ZN(new_n713_));
  INV_X1    g512(.A(G29gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n665_), .A2(new_n318_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(new_n351_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n653_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n479_), .A2(new_n714_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT106), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n713_), .A2(new_n714_), .B1(new_n717_), .B2(new_n719_), .ZN(G1328gat));
  OR2_X1    g519(.A1(new_n601_), .A2(KEYINPUT108), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n601_), .A2(KEYINPUT108), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n717_), .A2(G36gat), .A3(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT45), .Z(new_n726_));
  NAND3_X1  g525(.A1(new_n706_), .A2(new_n678_), .A3(new_n711_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n727_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT107), .B1(new_n727_), .B2(G36gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT46), .B(new_n726_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1329gat));
  INV_X1    g533(.A(G43gat), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n537_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n706_), .A2(new_n711_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n706_), .A2(KEYINPUT109), .A3(new_n711_), .A4(new_n736_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n717_), .B2(new_n537_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(G1330gat));
  NOR2_X1   g543(.A1(new_n717_), .A2(new_n446_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(G50gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n707_), .A2(new_n712_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n606_), .A2(G50gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(G1331gat));
  NOR2_X1   g548(.A1(new_n651_), .A2(new_n318_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n351_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n666_), .B2(new_n672_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G57gat), .B1(new_n753_), .B2(new_n611_), .ZN(new_n754_));
  NOR4_X1   g553(.A1(new_n320_), .A2(new_n635_), .A3(new_n651_), .A4(new_n660_), .ZN(new_n755_));
  INV_X1    g554(.A(G57gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n479_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1332gat));
  INV_X1    g557(.A(G64gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n723_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n752_), .A2(new_n723_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G64gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT48), .B(new_n759_), .C1(new_n752_), .C2(new_n723_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT111), .Z(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n752_), .B2(new_n603_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT49), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n755_), .A2(new_n767_), .A3(new_n603_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1334gat));
  INV_X1    g570(.A(G78gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n752_), .B2(new_n606_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT50), .Z(new_n774_));
  NAND2_X1  g573(.A1(new_n606_), .A2(new_n772_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT112), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n755_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(G1335gat));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n710_), .B(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n660_), .A2(new_n651_), .A3(new_n319_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782_), .B2(new_n611_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n635_), .A2(new_n651_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n660_), .A2(new_n715_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n786_), .A2(G85gat), .A3(new_n611_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n783_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT114), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n783_), .A2(new_n791_), .A3(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1336gat));
  OAI21_X1  g592(.A(G92gat), .B1(new_n782_), .B2(new_n724_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n601_), .A2(G92gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n784_), .A2(new_n785_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n794_), .A2(KEYINPUT115), .A3(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n782_), .B2(new_n537_), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n537_), .B(new_n786_), .C1(new_n203_), .C2(new_n204_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT51), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n802_), .A2(new_n807_), .A3(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1338gat));
  OR3_X1    g608(.A1(new_n786_), .A2(G106gat), .A3(new_n446_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n710_), .A2(new_n606_), .A3(new_n781_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G106gat), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(KEYINPUT52), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(KEYINPUT52), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n652_), .B2(new_n319_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n651_), .A2(new_n818_), .A3(new_n318_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NOR4_X1   g621(.A1(new_n702_), .A2(new_n820_), .A3(new_n351_), .A4(new_n822_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n351_), .A2(new_n819_), .A3(new_n817_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n821_), .B1(new_n824_), .B2(new_n291_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT12), .B1(new_n330_), .B2(new_n323_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n322_), .A2(new_n324_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT69), .B1(new_n830_), .B2(new_n327_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n326_), .A2(new_n321_), .A3(new_n328_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n827_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n328_), .A2(KEYINPUT118), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n328_), .A2(KEYINPUT55), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n326_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n326_), .B2(new_n834_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n833_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(KEYINPUT56), .A4(new_n343_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT55), .B1(new_n329_), .B2(new_n335_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n828_), .A2(new_n829_), .A3(new_n834_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n835_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n333_), .A2(new_n334_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n842_), .B1(new_n834_), .B2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT56), .B(new_n343_), .C1(new_n841_), .C2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT120), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n343_), .B1(new_n841_), .B2(new_n845_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n840_), .A2(new_n847_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n636_), .A2(new_n638_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n641_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n853_), .B2(new_n852_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n647_), .B1(new_n642_), .B2(new_n641_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n649_), .A2(new_n857_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n858_), .A2(new_n346_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n851_), .A2(KEYINPUT58), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n851_), .A2(new_n859_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n851_), .A2(KEYINPUT122), .A3(new_n859_), .A4(KEYINPUT58), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n862_), .A2(new_n865_), .A3(new_n702_), .A4(new_n866_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n347_), .A2(new_n858_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n651_), .A2(new_n346_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n850_), .B2(new_n846_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n289_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n872_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n867_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n826_), .B1(new_n875_), .B2(new_n318_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n446_), .A2(new_n601_), .A3(new_n479_), .A4(new_n603_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT59), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n867_), .A2(new_n874_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT124), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n867_), .A2(new_n881_), .A3(new_n874_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n873_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n826_), .B1(new_n883_), .B2(new_n318_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n877_), .A2(KEYINPUT123), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n877_), .A2(KEYINPUT123), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n885_), .A2(new_n886_), .A3(KEYINPUT59), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n651_), .B(new_n878_), .C1(new_n884_), .C2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G113gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n876_), .A2(new_n877_), .ZN(new_n890_));
  INV_X1    g689(.A(G113gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n651_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(G1340gat));
  OAI211_X1 g692(.A(new_n351_), .B(new_n878_), .C1(new_n884_), .C2(new_n887_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G120gat), .ZN(new_n895_));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n660_), .B2(KEYINPUT60), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n890_), .B(new_n897_), .C1(KEYINPUT60), .C2(new_n896_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(new_n898_), .ZN(G1341gat));
  OAI211_X1 g698(.A(new_n319_), .B(new_n878_), .C1(new_n884_), .C2(new_n887_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G127gat), .ZN(new_n901_));
  INV_X1    g700(.A(G127gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n890_), .A2(new_n902_), .A3(new_n319_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1342gat));
  OAI211_X1 g703(.A(new_n702_), .B(new_n878_), .C1(new_n884_), .C2(new_n887_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G134gat), .ZN(new_n906_));
  INV_X1    g705(.A(G134gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n890_), .A2(new_n907_), .A3(new_n665_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1343gat));
  NOR2_X1   g708(.A1(new_n876_), .A2(new_n446_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n723_), .A2(new_n611_), .A3(new_n603_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n651_), .A3(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n351_), .A3(new_n911_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n910_), .A2(new_n319_), .A3(new_n911_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n911_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G162gat), .B1(new_n919_), .B2(new_n291_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n289_), .A2(G162gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n919_), .B2(new_n921_), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n723_), .A2(new_n538_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n446_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n651_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G169gat), .B1(new_n884_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n826_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n867_), .A2(new_n881_), .A3(new_n874_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n881_), .B1(new_n867_), .B2(new_n874_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n873_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n931_), .B1(new_n935_), .B2(new_n319_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n936_), .A2(new_n559_), .A3(new_n651_), .A4(new_n926_), .ZN(new_n937_));
  OAI211_X1 g736(.A(KEYINPUT62), .B(G169gat), .C1(new_n884_), .C2(new_n927_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n930_), .A2(new_n937_), .A3(new_n938_), .ZN(G1348gat));
  OR2_X1    g738(.A1(new_n876_), .A2(new_n606_), .ZN(new_n940_));
  NOR4_X1   g739(.A1(new_n940_), .A2(new_n503_), .A3(new_n660_), .A4(new_n923_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n884_), .A2(new_n925_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n351_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n941_), .B1(new_n943_), .B2(new_n503_), .ZN(G1349gat));
  NOR2_X1   g743(.A1(new_n318_), .A2(new_n511_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n934_), .B1(new_n879_), .B2(KEYINPUT124), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n319_), .B1(new_n946_), .B2(new_n882_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n926_), .B(new_n945_), .C1(new_n947_), .C2(new_n826_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(KEYINPUT125), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n936_), .A2(new_n950_), .A3(new_n926_), .A4(new_n945_), .ZN(new_n951_));
  INV_X1    g750(.A(G183gat), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n924_), .A2(new_n319_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n940_), .B2(new_n953_), .ZN(new_n954_));
  AND3_X1   g753(.A1(new_n949_), .A2(new_n951_), .A3(new_n954_), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n936_), .A2(new_n702_), .A3(new_n926_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(G190gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n942_), .A2(new_n512_), .A3(new_n665_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1351gat));
  NOR3_X1   g758(.A1(new_n724_), .A2(new_n479_), .A3(new_n603_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n910_), .A2(new_n651_), .A3(new_n960_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g761(.A1(new_n910_), .A2(new_n351_), .A3(new_n960_), .ZN(new_n963_));
  XOR2_X1   g762(.A(KEYINPUT126), .B(G204gat), .Z(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1353gat));
  NOR2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(KEYINPUT127), .ZN(new_n967_));
  AND2_X1   g766(.A1(new_n910_), .A2(new_n960_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n318_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n967_), .B1(new_n968_), .B2(new_n969_), .ZN(new_n970_));
  AND4_X1   g769(.A1(new_n910_), .A2(new_n960_), .A3(new_n967_), .A4(new_n969_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n970_), .A2(new_n971_), .ZN(G1354gat));
  INV_X1    g771(.A(G218gat), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n968_), .A2(new_n973_), .A3(new_n665_), .ZN(new_n974_));
  AND3_X1   g773(.A1(new_n910_), .A2(new_n702_), .A3(new_n960_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n974_), .B1(new_n973_), .B2(new_n975_), .ZN(G1355gat));
endmodule


