//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_;
  NOR2_X1   g000(.A1(KEYINPUT69), .A2(G78gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT69), .A2(G78gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(G71gat), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G71gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(KEYINPUT69), .A2(G78gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(new_n202_), .ZN(new_n208_));
  INV_X1    g007(.A(G57gat), .ZN(new_n209_));
  INV_X1    g008(.A(G64gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G57gat), .A2(G64gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n205_), .A2(new_n208_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT70), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT70), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n205_), .A2(new_n208_), .A3(new_n214_), .A4(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n211_), .A2(new_n213_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(new_n212_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G99gat), .A2(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n235_), .A2(new_n226_), .A3(new_n236_), .A4(new_n237_), .ZN(new_n238_));
  AND3_X1   g037(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n233_), .B1(G99gat), .B2(G106gat), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n232_), .A2(new_n238_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G85gat), .B(G92gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT8), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n239_), .A2(new_n240_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT66), .B(KEYINPUT9), .Z(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G85gat), .A3(G92gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT10), .B(G99gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT65), .B1(new_n253_), .B2(G106gat), .ZN(new_n254_));
  OR3_X1    g053(.A1(new_n253_), .A2(KEYINPUT65), .A3(G106gat), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .A4(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n243_), .A2(KEYINPUT8), .A3(new_n244_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n247_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n225_), .A2(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n243_), .A2(KEYINPUT8), .A3(new_n244_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT8), .B1(new_n243_), .B2(new_n244_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n262_), .A2(new_n224_), .A3(new_n223_), .A4(new_n256_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n263_), .A3(KEYINPUT12), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT12), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n225_), .A2(new_n265_), .A3(new_n258_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(KEYINPUT64), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G120gat), .B(G148gat), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT5), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n270_), .A2(new_n272_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n269_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n282_), .B2(new_n271_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT13), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT83), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT22), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n277_), .A3(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT84), .Z(new_n294_));
  INV_X1    g093(.A(G183gat), .ZN(new_n295_));
  INV_X1    g094(.A(G190gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT23), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT85), .ZN(new_n298_));
  OR3_X1    g097(.A1(new_n295_), .A2(new_n296_), .A3(KEYINPUT23), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(KEYINPUT85), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(G183gat), .B2(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n294_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT82), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n289_), .A2(new_n277_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n310_), .B1(G169gat), .B2(G176gat), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n307_), .A2(KEYINPUT82), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n299_), .A2(new_n297_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n289_), .A3(new_n277_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n308_), .A2(new_n312_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n304_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT30), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G227gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT86), .ZN(new_n319_));
  XOR2_X1   g118(.A(G15gat), .B(G43gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G71gat), .B(G99gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n325_), .B(KEYINPUT87), .Z(new_n326_));
  NAND2_X1  g125(.A1(new_n317_), .A2(new_n324_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT88), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330_));
  INV_X1    g129(.A(G113gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G120gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n330_), .B(G113gat), .ZN(new_n334_));
  INV_X1    g133(.A(G120gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT31), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n329_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT3), .Z(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT2), .Z(new_n347_));
  OAI21_X1  g146(.A(new_n343_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT1), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n343_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n341_), .A2(KEYINPUT1), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n346_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n337_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n333_), .A2(new_n336_), .A3(new_n352_), .A4(new_n348_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT4), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(KEYINPUT4), .B2(new_n354_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT94), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n360_), .B2(new_n356_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT0), .B(G57gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(G85gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(G1gat), .B(G29gat), .Z(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(KEYINPUT99), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT99), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n362_), .A2(new_n372_), .A3(new_n369_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n340_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G211gat), .B(G218gat), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT21), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G197gat), .B(G204gat), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT90), .ZN(new_n381_));
  INV_X1    g180(.A(G197gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT89), .B1(new_n382_), .B2(G204gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(new_n378_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(new_n379_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n377_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n381_), .A2(new_n386_), .B1(KEYINPUT29), .B2(new_n353_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G50gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT28), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(G22gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n390_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n381_), .A2(new_n386_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n398_), .A2(new_n316_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n399_), .A2(KEYINPUT20), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n301_), .A2(new_n314_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT92), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT91), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n311_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n311_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n309_), .B1(new_n405_), .B2(KEYINPUT91), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n402_), .B(new_n307_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n313_), .B1(G183gat), .B2(G190gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT22), .B(G169gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n277_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n410_), .A3(new_n303_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n398_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT19), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n400_), .A2(new_n413_), .A3(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n412_), .A2(new_n398_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n398_), .A2(new_n316_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n418_), .A2(KEYINPUT20), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n417_), .B1(new_n420_), .B2(new_n416_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT18), .B(G64gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G92gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n418_), .A2(KEYINPUT20), .A3(new_n416_), .A4(new_n419_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n400_), .A2(new_n413_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n415_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n430_), .A3(new_n425_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(KEYINPUT27), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  INV_X1    g232(.A(new_n431_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n425_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n375_), .A2(new_n397_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n421_), .A2(KEYINPUT32), .A3(new_n425_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n428_), .A2(new_n430_), .A3(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n439_), .A2(new_n373_), .A3(new_n371_), .A4(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT95), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n370_), .A2(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n445_));
  NAND3_X1  g244(.A1(new_n362_), .A2(KEYINPUT95), .A3(new_n369_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n356_), .A2(KEYINPUT97), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n356_), .A2(KEYINPUT97), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n360_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n367_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT98), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n360_), .B2(new_n358_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n447_), .B(new_n453_), .C1(new_n454_), .C2(new_n370_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n435_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(KEYINPUT93), .A3(new_n431_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT93), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n442_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n374_), .A2(new_n397_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n461_), .A2(new_n397_), .B1(new_n462_), .B2(new_n437_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n438_), .B1(new_n463_), .B2(new_n339_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT73), .B(G29gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G36gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(G43gat), .B(G50gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n465_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT15), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G229gat), .A2(G233gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n468_), .A2(new_n472_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(new_n481_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n484_), .B(new_n481_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(G229gat), .A3(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G113gat), .B(G141gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G197gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT79), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(new_n289_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT80), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT81), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n464_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n225_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(new_n481_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n481_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G231gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G127gat), .B(G155gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(G183gat), .B(G211gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n509_), .B1(KEYINPUT17), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n514_), .B(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n518_), .B2(new_n509_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT34), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT75), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT75), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n525_), .B(new_n526_), .C1(new_n258_), .C2(new_n484_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n258_), .B2(new_n474_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n522_), .B(new_n523_), .C1(new_n527_), .C2(KEYINPUT74), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT76), .B(G134gat), .ZN(new_n531_));
  INV_X1    g330(.A(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(KEYINPUT36), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n528_), .A2(new_n529_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n530_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(KEYINPUT77), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(KEYINPUT36), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n536_), .B1(new_n530_), .B2(new_n537_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n541_), .B(new_n545_), .ZN(new_n546_));
  AND4_X1   g345(.A1(new_n287_), .A2(new_n503_), .A3(new_n520_), .A4(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n476_), .A3(new_n374_), .ZN(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n464_), .A2(new_n545_), .A3(new_n520_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n287_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n500_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT101), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT101), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n551_), .A2(new_n557_), .A3(new_n554_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n374_), .ZN(new_n560_));
  OAI21_X1  g359(.A(G1gat), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n550_), .A2(new_n561_), .ZN(G1324gat));
  OAI21_X1  g361(.A(G8gat), .B1(new_n555_), .B2(new_n437_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT39), .ZN(new_n564_));
  INV_X1    g363(.A(new_n437_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n547_), .A2(new_n477_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT40), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(G1325gat));
  OAI21_X1  g368(.A(G15gat), .B1(new_n559_), .B2(new_n340_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT41), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(G15gat), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n547_), .A2(new_n573_), .A3(new_n339_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(G1326gat));
  INV_X1    g374(.A(new_n397_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n547_), .A2(new_n394_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n578_), .B(G22gat), .C1(new_n559_), .C2(new_n397_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n397_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT102), .B1(new_n580_), .B2(new_n394_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n579_), .A2(KEYINPUT42), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT42), .B1(new_n579_), .B2(new_n581_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n577_), .B1(new_n582_), .B2(new_n583_), .ZN(G1327gat));
  XNOR2_X1  g383(.A(new_n541_), .B(new_n544_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT43), .B1(new_n546_), .B2(KEYINPUT103), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n464_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n464_), .B2(new_n585_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n554_), .B(new_n519_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT44), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n464_), .A2(new_n585_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n586_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n464_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n596_), .A2(KEYINPUT44), .A3(new_n554_), .A4(new_n519_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(G29gat), .A3(new_n374_), .ZN(new_n599_));
  INV_X1    g398(.A(G29gat), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n519_), .A2(new_n544_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT104), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n503_), .A2(new_n287_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n603_), .B2(new_n560_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n599_), .A2(new_n604_), .ZN(G1328gat));
  INV_X1    g404(.A(KEYINPUT107), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT106), .B1(new_n606_), .B2(KEYINPUT46), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n591_), .A2(new_n597_), .A3(new_n565_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G36gat), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n437_), .A2(G36gat), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n503_), .A2(new_n287_), .A3(new_n602_), .A4(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n607_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT106), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n609_), .A2(new_n615_), .A3(new_n613_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n606_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT46), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(G1329gat));
  NAND3_X1  g418(.A1(new_n598_), .A2(G43gat), .A3(new_n339_), .ZN(new_n620_));
  INV_X1    g419(.A(G43gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n603_), .B2(new_n340_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT108), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT47), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT47), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n620_), .A2(new_n626_), .A3(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(G1330gat));
  OR3_X1    g427(.A1(new_n603_), .A2(G50gat), .A3(new_n397_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n598_), .A2(new_n576_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT109), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(new_n631_), .A3(G50gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n630_), .B2(G50gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(G1331gat));
  NAND3_X1  g433(.A1(new_n551_), .A2(new_n552_), .A3(new_n501_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n635_), .A2(new_n209_), .A3(new_n560_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n464_), .A2(new_n553_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT110), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n552_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n546_), .A2(new_n520_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT111), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n639_), .A2(KEYINPUT111), .A3(new_n640_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n374_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n636_), .B1(new_n644_), .B2(new_n209_), .ZN(G1332gat));
  OAI21_X1  g444(.A(G64gat), .B1(new_n635_), .B2(new_n437_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT48), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n565_), .A2(new_n210_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n641_), .B2(new_n648_), .ZN(G1333gat));
  OAI21_X1  g448(.A(G71gat), .B1(new_n635_), .B2(new_n340_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT49), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n339_), .A2(new_n206_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n641_), .B2(new_n652_), .ZN(G1334gat));
  OAI21_X1  g452(.A(G78gat), .B1(new_n635_), .B2(new_n397_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT50), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n397_), .A2(G78gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n641_), .B2(new_n656_), .ZN(G1335gat));
  INV_X1    g456(.A(new_n639_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n602_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G85gat), .B1(new_n660_), .B2(new_n374_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n552_), .A2(new_n553_), .A3(new_n519_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT112), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT113), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n560_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n661_), .B1(new_n666_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g466(.A(G92gat), .B1(new_n660_), .B2(new_n565_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n665_), .A2(new_n437_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(G92gat), .ZN(G1337gat));
  NOR2_X1   g469(.A1(new_n340_), .A2(new_n253_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n660_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT51), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n227_), .B1(new_n664_), .B2(new_n339_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n672_), .A2(KEYINPUT114), .A3(new_n673_), .A4(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n671_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT114), .B1(new_n659_), .B2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT51), .B1(new_n678_), .B2(new_n674_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1338gat));
  NAND2_X1  g479(.A1(new_n576_), .A2(new_n228_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT52), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n664_), .A2(new_n576_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(G106gat), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT52), .B(new_n228_), .C1(new_n664_), .C2(new_n576_), .ZN(new_n685_));
  OAI22_X1  g484(.A1(new_n659_), .A2(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g486(.A(KEYINPUT119), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT118), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT55), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT115), .B1(new_n270_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT115), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n282_), .A2(new_n692_), .A3(KEYINPUT55), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n282_), .A2(KEYINPUT55), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n264_), .A2(new_n281_), .A3(new_n266_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n278_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n689_), .B1(new_n698_), .B2(KEYINPUT56), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n270_), .A2(KEYINPUT115), .A3(new_n690_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n692_), .B1(new_n282_), .B2(KEYINPUT55), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n695_), .A4(new_n696_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT117), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT117), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n702_), .A2(new_n705_), .A3(KEYINPUT56), .A4(new_n280_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT56), .B1(new_n702_), .B2(new_n280_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT118), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n699_), .A2(new_n704_), .A3(new_n706_), .A4(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n482_), .A2(new_n486_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(new_n483_), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n493_), .B(new_n711_), .C1(new_n483_), .C2(new_n488_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(new_n495_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n279_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT58), .B1(new_n709_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n688_), .B1(new_n716_), .B2(new_n546_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n704_), .A2(new_n706_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n702_), .A2(new_n280_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT56), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT118), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n689_), .B(KEYINPUT56), .C1(new_n702_), .C2(new_n280_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n714_), .B1(new_n718_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT58), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT119), .B(new_n585_), .C1(new_n724_), .C2(KEYINPUT58), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n717_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n286_), .A2(new_n713_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT116), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n703_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n500_), .B(new_n279_), .C1(new_n731_), .C2(new_n707_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n286_), .A2(KEYINPUT116), .A3(new_n713_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n734_), .A2(KEYINPUT57), .A3(new_n545_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT57), .B1(new_n734_), .B2(new_n545_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n727_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n519_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n501_), .A2(new_n546_), .A3(new_n287_), .A4(new_n520_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT54), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(KEYINPUT120), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT120), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n520_), .B1(new_n727_), .B2(new_n737_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n741_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n742_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n437_), .A2(new_n374_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(new_n340_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n397_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT59), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n576_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT59), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n749_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n751_), .A2(G113gat), .A3(new_n502_), .A4(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n331_), .B1(new_n750_), .B2(new_n553_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1340gat));
  INV_X1    g556(.A(new_n750_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n335_), .B1(new_n287_), .B2(KEYINPUT60), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n758_), .B(new_n759_), .C1(KEYINPUT60), .C2(new_n335_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n751_), .A2(new_n552_), .A3(new_n754_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n335_), .ZN(G1341gat));
  AOI21_X1  g561(.A(G127gat), .B1(new_n758_), .B2(new_n520_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n751_), .A2(new_n754_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n520_), .A2(G127gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT121), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n764_), .B2(new_n766_), .ZN(G1342gat));
  NAND4_X1  g566(.A1(new_n751_), .A2(G134gat), .A3(new_n585_), .A4(new_n754_), .ZN(new_n768_));
  INV_X1    g567(.A(G134gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n750_), .B2(new_n545_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1343gat));
  NOR2_X1   g570(.A1(new_n748_), .A2(new_n397_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n747_), .A2(new_n340_), .A3(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n553_), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n287_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g576(.A1(new_n773_), .A2(new_n519_), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT61), .B(G155gat), .Z(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1346gat));
  NOR3_X1   g579(.A1(new_n773_), .A2(new_n532_), .A3(new_n546_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n773_), .A2(new_n545_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n532_), .B2(new_n782_), .ZN(G1347gat));
  NAND2_X1  g582(.A1(new_n375_), .A2(new_n565_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT122), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n752_), .A2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n553_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(new_n289_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n788_), .A2(KEYINPUT62), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n409_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(KEYINPUT62), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(new_n790_), .A3(new_n791_), .ZN(G1348gat));
  INV_X1    g591(.A(new_n786_), .ZN(new_n793_));
  AOI21_X1  g592(.A(G176gat), .B1(new_n793_), .B2(new_n552_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n742_), .A2(new_n397_), .A3(new_n746_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT123), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT123), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n742_), .A2(new_n746_), .A3(new_n797_), .A4(new_n397_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n799_), .A2(G176gat), .A3(new_n785_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n794_), .B1(new_n800_), .B2(new_n552_), .ZN(G1349gat));
  NOR3_X1   g600(.A1(new_n786_), .A2(new_n305_), .A3(new_n519_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n785_), .A2(new_n520_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT124), .B1(new_n799_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n806_), .B(new_n803_), .C1(new_n796_), .C2(new_n798_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n802_), .B1(new_n808_), .B2(new_n295_), .ZN(G1350gat));
  OAI21_X1  g608(.A(G190gat), .B1(new_n786_), .B2(new_n546_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n544_), .A2(new_n306_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n786_), .B2(new_n811_), .ZN(G1351gat));
  NOR3_X1   g611(.A1(new_n437_), .A2(new_n374_), .A3(new_n397_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n742_), .A2(new_n746_), .A3(new_n340_), .A4(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n553_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT126), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT126), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT125), .B(new_n818_), .C1(new_n814_), .C2(new_n553_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n816_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n382_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n817_), .A2(new_n821_), .A3(new_n382_), .A4(new_n819_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1352gat));
  NOR2_X1   g624(.A1(new_n814_), .A2(new_n287_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(new_n274_), .ZN(G1353gat));
  INV_X1    g626(.A(new_n814_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n520_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n830_));
  AND2_X1   g629(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n829_), .B2(new_n830_), .ZN(G1354gat));
  AOI21_X1  g632(.A(G218gat), .B1(new_n828_), .B2(new_n544_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n585_), .A2(G218gat), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT127), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n828_), .B2(new_n836_), .ZN(G1355gat));
endmodule


