//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n204_));
  INV_X1    g003(.A(G85gat), .ZN(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  OAI211_X1 g006(.A(G85gat), .B(G92gat), .C1(KEYINPUT66), .C2(KEYINPUT9), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n203_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n207_), .A2(new_n208_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT10), .B(G99gat), .Z(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT65), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n212_), .A2(KEYINPUT65), .A3(new_n213_), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n210_), .B(new_n211_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  OR3_X1    g017(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n203_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G85gat), .B(G92gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT67), .ZN(new_n222_));
  AND4_X1   g021(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  AOI22_X1  g022(.A1(new_n220_), .A2(new_n221_), .B1(new_n222_), .B2(new_n217_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n216_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT68), .B(G71gat), .Z(new_n226_));
  INV_X1    g025(.A(G78gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(G71gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G78gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n228_), .A2(new_n230_), .B1(KEYINPUT11), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(KEYINPUT11), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n229_), .B(new_n227_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n225_), .A2(new_n236_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n235_), .B(new_n216_), .C1(new_n224_), .C2(new_n223_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT12), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n225_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G230gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT64), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G120gat), .B(G148gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT5), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G176gat), .B(G204gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n245_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n244_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n254_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(new_n246_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n253_), .A2(KEYINPUT69), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT69), .B1(new_n253_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT13), .ZN(new_n260_));
  XOR2_X1   g059(.A(G8gat), .B(G36gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(G64gat), .B(G92gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n266_));
  AND2_X1   g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT22), .B(G169gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT90), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT90), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT22), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(G169gat), .ZN(new_n273_));
  INV_X1    g072(.A(G169gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT22), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G183gat), .ZN(new_n282_));
  INV_X1    g081(.A(G190gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n281_), .A2(new_n284_), .B1(G169gat), .B2(G176gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n278_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT25), .B(G183gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT26), .B(G190gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT24), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(G169gat), .B2(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n274_), .A2(new_n277_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n286_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G197gat), .A2(G204gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G197gat), .A2(G204gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(KEYINPUT21), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT21), .ZN(new_n306_));
  INV_X1    g105(.A(new_n304_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n302_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G211gat), .B(G218gat), .Z(new_n311_));
  NAND4_X1  g110(.A1(new_n311_), .A2(KEYINPUT21), .A3(new_n303_), .A4(new_n304_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT20), .B1(new_n301_), .B2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n310_), .A2(new_n312_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n269_), .A2(KEYINPUT83), .A3(new_n277_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT83), .B1(new_n269_), .B2(new_n277_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n285_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n282_), .A2(KEYINPUT25), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT25), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G183gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n283_), .A2(KEYINPUT26), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G190gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT82), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT82), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n327_), .A2(new_n281_), .A3(new_n299_), .A4(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n315_), .B1(new_n318_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n268_), .B1(new_n314_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n301_), .B2(new_n313_), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n268_), .B(KEYINPUT89), .Z(new_n334_));
  NAND3_X1  g133(.A1(new_n315_), .A2(new_n318_), .A3(new_n329_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n265_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT94), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n268_), .B(KEYINPUT89), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n278_), .A2(new_n285_), .B1(new_n294_), .B2(new_n299_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT20), .B1(new_n341_), .B2(new_n315_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n315_), .A2(new_n318_), .A3(new_n329_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n340_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n332_), .B1(new_n341_), .B2(new_n315_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n318_), .A2(new_n329_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n313_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n268_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n349_), .A3(new_n265_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n338_), .A2(new_n339_), .A3(KEYINPUT27), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(KEYINPUT27), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT94), .B1(new_n352_), .B2(new_n337_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n265_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n357_), .B2(new_n350_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G22gat), .B(G50gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT28), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT1), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT85), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370_));
  NAND3_X1  g169(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n366_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT84), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(G141gat), .A3(G148gat), .ZN(new_n379_));
  INV_X1    g178(.A(G141gat), .ZN(new_n380_));
  INV_X1    g179(.A(G148gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n375_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n373_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT2), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n377_), .A2(new_n379_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n386_), .B1(new_n388_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n385_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n385_), .B2(new_n394_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n363_), .B1(new_n398_), .B2(KEYINPUT29), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n362_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(KEYINPUT87), .A3(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G78gat), .B(G106gat), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n399_), .A2(KEYINPUT87), .A3(new_n401_), .A4(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n399_), .A2(new_n401_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n398_), .A2(KEYINPUT29), .ZN(new_n411_));
  AND2_X1   g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n315_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n369_), .A2(new_n371_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n373_), .B1(new_n414_), .B2(KEYINPUT1), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n383_), .B1(new_n415_), .B2(new_n372_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n374_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n377_), .A2(new_n379_), .A3(new_n387_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT29), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n313_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n411_), .A2(new_n413_), .B1(new_n412_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n410_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n407_), .A2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n404_), .A2(new_n410_), .A3(new_n423_), .A4(new_n406_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n360_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G43gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n346_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G127gat), .B(G134gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G113gat), .B(G120gat), .Z(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G113gat), .B(G120gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n431_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n431_), .A2(new_n438_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(G15gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT30), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT31), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OR3_X1    g245(.A1(new_n439_), .A2(new_n440_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n385_), .A2(new_n394_), .A3(new_n438_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n385_), .A2(new_n438_), .A3(new_n394_), .A4(KEYINPUT92), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT86), .B1(new_n416_), .B2(new_n420_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n385_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n438_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n454_), .A2(KEYINPUT4), .A3(new_n458_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT4), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n455_), .A2(new_n462_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n459_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n460_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G1gat), .B(G29gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G85gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT0), .B(G57gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n460_), .B(new_n470_), .C1(new_n461_), .C2(new_n465_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n449_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n428_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n473_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n463_), .A2(new_n464_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n454_), .A2(new_n458_), .A3(KEYINPUT4), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n470_), .B1(new_n480_), .B2(new_n460_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n265_), .A2(KEYINPUT32), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n344_), .A2(new_n349_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n331_), .A2(new_n336_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n483_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT93), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n488_));
  AOI211_X1 g287(.A(new_n488_), .B(new_n483_), .C1(new_n331_), .C2(new_n336_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n484_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n344_), .A2(new_n349_), .A3(new_n265_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(new_n356_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n470_), .A2(KEYINPUT33), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n460_), .B(new_n493_), .C1(new_n461_), .C2(new_n465_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n454_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n463_), .A2(new_n459_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n471_), .B(new_n495_), .C1(new_n461_), .C2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n398_), .A2(new_n457_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n479_), .A2(new_n478_), .B1(new_n499_), .B2(new_n459_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT33), .B1(new_n500_), .B2(new_n470_), .ZN(new_n501_));
  OAI22_X1  g300(.A1(new_n482_), .A2(new_n490_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n426_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n404_), .A2(new_n406_), .B1(new_n410_), .B2(new_n423_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n474_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n358_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n502_), .A2(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n449_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n476_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT34), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT35), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT70), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n513_), .A2(KEYINPUT35), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(KEYINPUT73), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(KEYINPUT73), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G29gat), .B(G36gat), .Z(new_n520_));
  INV_X1    g319(.A(KEYINPUT71), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G29gat), .B(G36gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT71), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI221_X1 g328(.A(new_n519_), .B1(new_n511_), .B2(new_n515_), .C1(new_n225_), .C2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n522_), .A2(new_n524_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n525_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n225_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n511_), .B(new_n515_), .C1(new_n530_), .C2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n225_), .A2(new_n529_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n519_), .B1(new_n515_), .B2(new_n511_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n515_), .A2(new_n511_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n539_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G190gat), .B(G218gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT74), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n547_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n551_), .B(KEYINPUT36), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n541_), .A2(new_n546_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT37), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n557_), .B2(KEYINPUT76), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n555_), .B(new_n557_), .C1(KEYINPUT76), .C2(new_n559_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564_));
  INV_X1    g363(.A(G1gat), .ZN(new_n565_));
  INV_X1    g364(.A(G8gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT14), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G1gat), .B(G8gat), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n569_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT77), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n235_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  XOR2_X1   g376(.A(G127gat), .B(G155gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT16), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n576_), .A2(new_n577_), .A3(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(KEYINPUT17), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n563_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT81), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G169gat), .B(G197gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  NAND3_X1  g389(.A1(new_n528_), .A2(new_n571_), .A3(new_n570_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT80), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n538_), .A2(new_n536_), .A3(new_n572_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT79), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n538_), .A2(new_n536_), .A3(KEYINPUT79), .A4(new_n572_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n572_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n572_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n533_), .A2(new_n534_), .B1(new_n571_), .B2(new_n570_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT78), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n592_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n590_), .B1(new_n600_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n590_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n599_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n587_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n600_), .A2(new_n608_), .A3(new_n590_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n599_), .B2(new_n607_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(KEYINPUT81), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n260_), .A2(new_n510_), .A3(new_n586_), .A4(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n620_), .A2(new_n565_), .A3(new_n474_), .A4(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n260_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n625_), .A2(new_n616_), .A3(new_n585_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n505_), .A2(new_n507_), .A3(new_n475_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n502_), .A2(new_n505_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n427_), .A2(new_n507_), .A3(new_n482_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n627_), .B1(new_n630_), .B2(new_n449_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n558_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n565_), .B1(new_n635_), .B2(new_n474_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n624_), .A2(new_n636_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n622_), .A2(KEYINPUT97), .A3(new_n623_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT97), .B1(new_n622_), .B2(new_n623_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(G1324gat));
  NAND4_X1  g441(.A1(new_n620_), .A2(new_n566_), .A3(new_n360_), .A4(new_n621_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT99), .Z(new_n644_));
  OAI21_X1  g443(.A(G8gat), .B1(new_n634_), .B2(new_n507_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT39), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n634_), .B2(new_n449_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT41), .Z(new_n651_));
  AND2_X1   g450(.A1(new_n620_), .A2(new_n621_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n442_), .A3(new_n509_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(KEYINPUT100), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(KEYINPUT100), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n654_), .A3(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n635_), .B2(new_n427_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(KEYINPUT42), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n652_), .A2(new_n657_), .A3(new_n427_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT42), .B1(new_n660_), .B2(new_n661_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n585_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n558_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n260_), .A2(new_n510_), .A3(new_n617_), .A4(new_n668_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n669_), .A2(KEYINPUT104), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(KEYINPUT104), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G29gat), .B1(new_n672_), .B2(new_n474_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n509_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n674_), .B(new_n563_), .C1(new_n675_), .C2(new_n627_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT102), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n510_), .A2(new_n678_), .A3(new_n674_), .A4(new_n563_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n563_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT43), .B1(new_n631_), .B2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n677_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n625_), .A2(new_n616_), .A3(new_n667_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT103), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n682_), .A2(new_n686_), .A3(KEYINPUT44), .A4(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n682_), .A2(new_n683_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n688_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n474_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n673_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  INV_X1    g494(.A(G36gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n507_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n688_), .B2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n670_), .A2(new_n696_), .A3(new_n360_), .A4(new_n671_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n695_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n695_), .B(KEYINPUT46), .C1(new_n698_), .C2(new_n701_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  AND4_X1   g505(.A1(G43gat), .A2(new_n688_), .A3(new_n509_), .A4(new_n691_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n670_), .A2(new_n509_), .A3(new_n671_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT106), .B(G43gat), .Z(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT107), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OR3_X1    g512(.A1(new_n707_), .A2(new_n711_), .A3(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n707_), .B2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n672_), .B2(new_n427_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n427_), .A2(G50gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n692_), .B2(new_n718_), .ZN(G1331gat));
  NAND3_X1  g518(.A1(new_n625_), .A2(new_n510_), .A3(new_n616_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n563_), .A3(new_n585_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n474_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n260_), .A2(new_n617_), .A3(new_n585_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n633_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n482_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1332gat));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n721_), .A2(new_n728_), .A3(new_n360_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G64gat), .B1(new_n725_), .B2(new_n507_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT48), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT48), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(new_n732_), .ZN(G1333gat));
  NOR2_X1   g532(.A1(new_n449_), .A2(G71gat), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT109), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n721_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G71gat), .B1(new_n725_), .B2(new_n449_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(KEYINPUT49), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(KEYINPUT49), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(G1334gat));
  NAND3_X1  g539(.A1(new_n721_), .A2(new_n227_), .A3(new_n427_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n724_), .A2(new_n427_), .A3(new_n633_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(G78gat), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G78gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1335gat));
  NOR3_X1   g545(.A1(new_n720_), .A2(new_n558_), .A3(new_n667_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n205_), .A3(new_n474_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n260_), .A2(new_n617_), .A3(new_n667_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n682_), .A2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n474_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n751_), .B2(new_n205_), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n747_), .A2(new_n206_), .A3(new_n360_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n750_), .A2(new_n360_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n206_), .ZN(G1337gat));
  NAND2_X1  g554(.A1(new_n750_), .A2(new_n509_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n509_), .A2(new_n212_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n756_), .A2(G99gat), .B1(new_n747_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(KEYINPUT113), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT113), .B1(new_n758_), .B2(new_n759_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n758_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT51), .B1(new_n758_), .B2(new_n762_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n760_), .A2(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n747_), .A2(new_n213_), .A3(new_n427_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n682_), .A2(KEYINPUT114), .A3(new_n427_), .A4(new_n749_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(G106gat), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n682_), .A2(new_n427_), .A3(new_n749_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n768_), .A2(new_n769_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n769_), .B1(new_n768_), .B2(new_n772_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n766_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT53), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n766_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1339gat));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n428_), .A2(new_n474_), .A3(new_n509_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n260_), .A2(new_n586_), .A3(new_n616_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n612_), .A2(new_n615_), .A3(new_n253_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n239_), .A2(new_n254_), .A3(new_n241_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n255_), .B1(KEYINPUT55), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n242_), .A2(KEYINPUT55), .A3(new_n244_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n251_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT56), .B(new_n251_), .C1(new_n788_), .C2(new_n790_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n786_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n604_), .B(new_n593_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n603_), .A2(new_n606_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n593_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n610_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n613_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n257_), .A2(new_n258_), .A3(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n558_), .B1(new_n795_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n558_), .B(new_n803_), .C1(new_n795_), .C2(new_n801_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n794_), .A2(KEYINPUT117), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n787_), .A2(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n245_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n789_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(KEYINPUT56), .A4(new_n251_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n808_), .A2(new_n813_), .A3(new_n793_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n255_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n800_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n814_), .A2(KEYINPUT58), .A3(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n563_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n667_), .B1(new_n807_), .B2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n780_), .B(new_n782_), .C1(new_n785_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n820_), .A2(new_n563_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n818_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n824_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n819_), .A2(KEYINPUT119), .A3(new_n563_), .A4(new_n820_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n807_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n585_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n784_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n783_), .B(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n781_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n823_), .B1(new_n834_), .B2(new_n780_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n616_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n834_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n616_), .A2(G113gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1340gat));
  OAI211_X1 g638(.A(new_n625_), .B(new_n823_), .C1(new_n834_), .C2(new_n780_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G120gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n260_), .A2(KEYINPUT60), .ZN(new_n842_));
  MUX2_X1   g641(.A(new_n842_), .B(KEYINPUT60), .S(G120gat), .Z(new_n843_));
  AOI22_X1  g642(.A1(new_n821_), .A2(new_n824_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n667_), .B1(new_n844_), .B2(new_n829_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n782_), .B(new_n843_), .C1(new_n845_), .C2(new_n785_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n834_), .A2(KEYINPUT120), .A3(new_n843_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n841_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n841_), .A2(new_n850_), .A3(KEYINPUT121), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n835_), .B2(new_n585_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n585_), .A2(G127gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n837_), .B2(new_n857_), .ZN(G1342gat));
  OAI21_X1  g657(.A(G134gat), .B1(new_n835_), .B2(new_n680_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n558_), .A2(G134gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n837_), .B2(new_n860_), .ZN(G1343gat));
  NOR4_X1   g660(.A1(new_n505_), .A2(new_n360_), .A3(new_n482_), .A4(new_n509_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n845_), .B2(new_n785_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n616_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(new_n380_), .ZN(G1344gat));
  NOR2_X1   g664(.A1(new_n863_), .A2(new_n260_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(new_n381_), .ZN(G1345gat));
  NOR2_X1   g666(.A1(new_n863_), .A2(new_n585_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT61), .B(G155gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1346gat));
  OAI21_X1  g669(.A(G162gat), .B1(new_n863_), .B2(new_n680_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n558_), .A2(G162gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n863_), .B2(new_n872_), .ZN(G1347gat));
  OR2_X1    g672(.A1(new_n785_), .A2(new_n822_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n360_), .A2(new_n475_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n427_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT122), .B1(new_n877_), .B2(new_n616_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n874_), .A2(new_n879_), .A3(new_n617_), .A4(new_n876_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(G169gat), .A3(new_n880_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n877_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n884_), .A2(new_n276_), .A3(new_n270_), .A4(new_n617_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n882_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n878_), .A2(G169gat), .A3(new_n886_), .A4(new_n880_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n883_), .A2(new_n885_), .A3(new_n887_), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n884_), .B2(new_n625_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n845_), .A2(new_n785_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n427_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n260_), .A2(new_n277_), .A3(new_n875_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n891_), .B2(new_n892_), .ZN(G1349gat));
  NOR3_X1   g692(.A1(new_n877_), .A2(new_n292_), .A3(new_n585_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n891_), .A2(new_n360_), .A3(new_n475_), .A4(new_n667_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n282_), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n877_), .B2(new_n680_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n632_), .A2(new_n293_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT124), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n877_), .B2(new_n899_), .ZN(G1351gat));
  NAND3_X1  g699(.A1(new_n506_), .A2(new_n360_), .A3(new_n449_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n890_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n617_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n625_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g705(.A(new_n585_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n907_));
  OR2_X1    g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n902_), .A2(new_n907_), .B1(KEYINPUT125), .B2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(KEYINPUT125), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT126), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n909_), .B(new_n911_), .ZN(G1354gat));
  AOI21_X1  g711(.A(G218gat), .B1(new_n902_), .B2(new_n632_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n563_), .A2(G218gat), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT127), .Z(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n902_), .B2(new_n915_), .ZN(G1355gat));
endmodule


