//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT92), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT91), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n204_), .B1(new_n205_), .B2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(new_n205_), .B2(new_n210_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n206_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n213_), .A2(new_n214_), .A3(new_n208_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(KEYINPUT1), .B2(new_n202_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G113gat), .B(G120gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT90), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n219_), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n225_), .A2(KEYINPUT4), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT102), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n223_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n212_), .A2(new_n216_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(KEYINPUT4), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n226_), .B1(new_n227_), .B2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n225_), .A2(new_n229_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(KEYINPUT102), .A3(KEYINPUT4), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT103), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G1gat), .B(G29gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT0), .ZN(new_n239_));
  INV_X1    g038(.A(G57gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G85gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n232_), .A2(new_n236_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n243_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n236_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n249_), .B2(new_n244_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G8gat), .B(G36gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT18), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G64gat), .ZN(new_n254_));
  INV_X1    g053(.A(G92gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT25), .B(G183gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT84), .ZN(new_n261_));
  INV_X1    g060(.A(G169gat), .ZN(new_n262_));
  INV_X1    g061(.A(G176gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(KEYINPUT24), .A3(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n264_), .A2(KEYINPUT24), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT23), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n261_), .A2(new_n266_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT86), .B(G176gat), .Z(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT85), .B1(new_n262_), .B2(KEYINPUT22), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT22), .B(G169gat), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n271_), .B(new_n272_), .C1(KEYINPUT85), .C2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT87), .B1(new_n268_), .B2(KEYINPUT23), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n269_), .B2(KEYINPUT87), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n265_), .B(new_n274_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n270_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n270_), .A2(KEYINPUT88), .A3(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G204gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT95), .B1(new_n284_), .B2(G197gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT95), .ZN(new_n286_));
  INV_X1    g085(.A(G197gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(G204gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n285_), .B(new_n288_), .C1(new_n287_), .C2(G204gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT98), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G211gat), .B(G218gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT97), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT21), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n292_), .B2(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n284_), .A2(G197gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n287_), .A2(G204gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT21), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n298_), .B(new_n291_), .C1(new_n289_), .C2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n283_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G226gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT19), .ZN(new_n304_));
  INV_X1    g103(.A(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n271_), .A2(new_n273_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n269_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n265_), .B(new_n306_), .C1(new_n307_), .C2(new_n277_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n310_), .B(new_n260_), .C1(new_n264_), .C2(new_n309_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n311_), .B2(new_n276_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT20), .B1(new_n305_), .B2(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n302_), .A2(new_n304_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n304_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n283_), .A2(new_n301_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n305_), .B2(new_n313_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n257_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n304_), .B1(new_n302_), .B2(new_n314_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n256_), .A3(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n321_), .A2(KEYINPUT27), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT105), .B(KEYINPUT27), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n257_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n327_), .B1(new_n329_), .B2(new_n324_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n251_), .A2(new_n325_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n224_), .B(KEYINPUT31), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G71gat), .B(G99gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G15gat), .B(G43gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n281_), .A2(KEYINPUT30), .A3(new_n282_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT30), .B1(new_n281_), .B2(new_n282_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n337_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n283_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n338_), .A3(new_n336_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT89), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(new_n344_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n335_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n341_), .A2(new_n344_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n346_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n334_), .A3(new_n348_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n217_), .A2(KEYINPUT29), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n356_), .A2(KEYINPUT94), .A3(new_n357_), .A4(new_n301_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n301_), .A2(KEYINPUT94), .ZN(new_n361_));
  OAI211_X1 g160(.A(G228gat), .B(G233gat), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n358_), .B2(new_n362_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT100), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n364_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT99), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n212_), .A2(new_n359_), .A3(new_n216_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n375_));
  XNOR2_X1  g174(.A(G22gat), .B(G50gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n374_), .B(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n370_), .B1(new_n373_), .B2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n378_), .B(new_n370_), .C1(new_n367_), .C2(KEYINPUT99), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n369_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n367_), .A2(KEYINPUT99), .ZN(new_n383_));
  INV_X1    g182(.A(new_n378_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT100), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n368_), .A3(new_n380_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n355_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n355_), .B1(new_n386_), .B2(new_n382_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n331_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n250_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n324_), .A3(new_n329_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n247_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n250_), .B2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n246_), .A2(new_n250_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n256_), .A2(KEYINPUT32), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n322_), .A2(new_n323_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT104), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(KEYINPUT32), .B(new_n256_), .C1(new_n315_), .C2(new_n320_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n399_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n392_), .A2(new_n395_), .B1(new_n396_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n382_), .A2(new_n386_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n405_), .A2(new_n355_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n389_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT17), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G127gat), .B(G155gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT16), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G183gat), .ZN(new_n412_));
  INV_X1    g211(.A(G211gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G1gat), .ZN(new_n415_));
  INV_X1    g214(.A(G8gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT14), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n417_), .A2(KEYINPUT79), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G15gat), .B(G22gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(KEYINPUT79), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G1gat), .B(G8gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G71gat), .B(G78gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G57gat), .B(G64gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT11), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(KEYINPUT11), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n423_), .B(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(G231gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI211_X1 g233(.A(new_n409_), .B(new_n414_), .C1(new_n434_), .C2(KEYINPUT80), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(KEYINPUT80), .B2(new_n434_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n414_), .B(KEYINPUT17), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT81), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n242_), .A2(new_n255_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n445_));
  INV_X1    g244(.A(G99gat), .ZN(new_n446_));
  INV_X1    g245(.A(G106gat), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .A4(KEYINPUT67), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  OAI22_X1  g248(.A1(new_n449_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G99gat), .A2(G106gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n444_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT8), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT69), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT69), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n460_), .A3(KEYINPUT8), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n448_), .A2(new_n450_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n444_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT68), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT68), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n462_), .A2(new_n466_), .A3(new_n463_), .A4(new_n444_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n459_), .A2(new_n461_), .A3(new_n465_), .A4(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n456_), .B1(new_n474_), .B2(new_n447_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT9), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n442_), .A2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT66), .B(new_n477_), .C1(new_n444_), .C2(new_n476_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n476_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n477_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n475_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G29gat), .B(G36gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G43gat), .B(G50gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n468_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n465_), .A2(new_n467_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n460_), .B1(new_n457_), .B2(KEYINPUT8), .ZN(new_n491_));
  AOI211_X1 g290(.A(KEYINPUT69), .B(new_n463_), .C1(new_n462_), .C2(new_n444_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n490_), .A2(new_n493_), .B1(new_n483_), .B2(new_n475_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n487_), .B(KEYINPUT15), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n489_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT75), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G232gat), .A2(G233gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT34), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n468_), .A2(new_n484_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n495_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n500_), .B(new_n502_), .C1(new_n505_), .C2(new_n489_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n502_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n496_), .B2(KEYINPUT75), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n499_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n468_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n495_), .B1(new_n468_), .B2(new_n484_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT75), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n502_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n496_), .A2(KEYINPUT75), .A3(new_n507_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(KEYINPUT35), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT77), .B1(new_n509_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n506_), .A2(new_n508_), .A3(new_n497_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n498_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT36), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G190gat), .B(G218gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT76), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(G134gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G162gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n517_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n524_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n509_), .A2(new_n515_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n531_), .B2(KEYINPUT36), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n532_), .A2(new_n516_), .A3(new_n527_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT37), .B1(new_n529_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n525_), .A2(new_n517_), .A3(new_n528_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n516_), .B1(new_n532_), .B2(new_n527_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT78), .B(KEYINPUT37), .Z(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n408_), .A2(new_n440_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n494_), .A2(new_n430_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n430_), .B1(new_n468_), .B2(new_n484_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n430_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n503_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n550_));
  AOI211_X1 g349(.A(new_n430_), .B(new_n550_), .C1(new_n468_), .C2(new_n484_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n541_), .B(new_n549_), .C1(new_n551_), .C2(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT64), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  MUX2_X1   g354(.A(new_n544_), .B(new_n552_), .S(new_n555_), .Z(new_n556_));
  XNOR2_X1  g355(.A(G120gat), .B(G148gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT72), .ZN(new_n558_));
  XOR2_X1   g357(.A(G176gat), .B(G204gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n556_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n556_), .A2(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n564_), .B(new_n565_), .C1(KEYINPUT73), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(KEYINPUT74), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT74), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n504_), .A2(new_n423_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n423_), .A2(new_n487_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n423_), .B(new_n487_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT82), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G169gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n287_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT83), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n585_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n575_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n540_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n396_), .B(KEYINPUT106), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n415_), .A3(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n535_), .A2(new_n536_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n389_), .B2(new_n407_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT109), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n591_), .B(new_n440_), .C1(new_n572_), .C2(new_n574_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT108), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n396_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n595_), .A2(new_n596_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  NOR2_X1   g406(.A1(new_n325_), .A2(new_n330_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n593_), .A2(new_n416_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(new_n609_), .A3(new_n603_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n611_), .A2(new_n612_), .A3(G8gat), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n611_), .B2(G8gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT40), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(G1325gat));
  INV_X1    g416(.A(G15gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n593_), .A2(new_n618_), .A3(new_n355_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n601_), .A2(new_n355_), .A3(new_n603_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n620_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT41), .B1(new_n620_), .B2(G15gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n619_), .B1(new_n621_), .B2(new_n622_), .ZN(G1326gat));
  INV_X1    g422(.A(G22gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n593_), .A2(new_n624_), .A3(new_n405_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n405_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G22gat), .B1(new_n604_), .B2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(KEYINPUT42), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(KEYINPUT42), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n625_), .B1(new_n628_), .B2(new_n629_), .ZN(G1327gat));
  NOR2_X1   g429(.A1(new_n592_), .A2(new_n440_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n598_), .B1(new_n389_), .B2(new_n407_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n251_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  INV_X1    g435(.A(new_n539_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n408_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT110), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n408_), .A2(KEYINPUT110), .A3(new_n636_), .A4(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n408_), .A2(new_n637_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT43), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n640_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n631_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(G29gat), .A3(new_n594_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT44), .B1(new_n644_), .B2(new_n631_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n635_), .B1(new_n646_), .B2(new_n648_), .ZN(G1328gat));
  XNOR2_X1  g448(.A(new_n608_), .B(KEYINPUT111), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  OR3_X1    g450(.A1(new_n633_), .A2(KEYINPUT45), .A3(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT45), .B1(new_n633_), .B2(new_n651_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n652_), .A2(new_n653_), .B1(KEYINPUT112), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n645_), .A2(new_n609_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G36gat), .B1(new_n656_), .B2(new_n647_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n654_), .A2(KEYINPUT112), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n655_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1329gat));
  NAND3_X1  g460(.A1(new_n645_), .A2(G43gat), .A3(new_n355_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n355_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n633_), .A2(new_n663_), .ZN(new_n664_));
  OAI22_X1  g463(.A1(new_n662_), .A2(new_n647_), .B1(G43gat), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g465(.A(G50gat), .B1(new_n634_), .B2(new_n405_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n645_), .A2(G50gat), .A3(new_n405_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(new_n648_), .ZN(G1331gat));
  INV_X1    g468(.A(new_n440_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n575_), .A2(new_n591_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n601_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G57gat), .B1(new_n672_), .B2(new_n396_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n540_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n575_), .A2(new_n591_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n594_), .A2(new_n240_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1332gat));
  OAI21_X1  g477(.A(G64gat), .B1(new_n672_), .B2(new_n650_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT48), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n650_), .A2(G64gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n676_), .B2(new_n681_), .ZN(G1333gat));
  OAI21_X1  g481(.A(G71gat), .B1(new_n672_), .B2(new_n663_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT49), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n663_), .A2(G71gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n676_), .B2(new_n685_), .ZN(G1334gat));
  OAI21_X1  g485(.A(G78gat), .B1(new_n672_), .B2(new_n626_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT50), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n626_), .A2(G78gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n676_), .B2(new_n689_), .ZN(G1335gat));
  NOR3_X1   g489(.A1(new_n575_), .A2(new_n591_), .A3(new_n440_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n632_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n594_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n242_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT113), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n644_), .A2(new_n691_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT114), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n396_), .A2(new_n242_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(G1336gat));
  INV_X1    g499(.A(new_n692_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n255_), .A3(new_n609_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n650_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n698_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n704_), .B2(new_n255_), .ZN(G1337gat));
  NAND3_X1  g504(.A1(new_n701_), .A2(new_n474_), .A3(new_n355_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n644_), .A2(new_n355_), .A3(new_n691_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT115), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G99gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G99gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT51), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n706_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1338gat));
  NAND3_X1  g514(.A1(new_n701_), .A2(new_n447_), .A3(new_n405_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n644_), .A2(new_n405_), .A3(new_n691_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(G106gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n717_), .B2(G106gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT53), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT53), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n723_), .B(new_n716_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1339gat));
  NAND2_X1  g524(.A1(new_n591_), .A2(new_n565_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT116), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n549_), .A2(new_n541_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n550_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n548_), .B1(new_n543_), .B2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n727_), .B(new_n554_), .C1(new_n728_), .C2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n727_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n728_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n730_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(KEYINPUT55), .A4(new_n555_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n562_), .B1(new_n734_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT56), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n736_), .B(new_n739_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n562_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n726_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n583_), .A2(new_n588_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n576_), .A2(new_n577_), .A3(new_n581_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n580_), .A2(new_n578_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n588_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT57), .B(new_n598_), .C1(new_n746_), .C2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT120), .ZN(new_n754_));
  INV_X1    g553(.A(new_n752_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n562_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n562_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n758_), .B2(new_n726_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(KEYINPUT57), .A4(new_n598_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n754_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n751_), .B1(new_n556_), .B2(new_n563_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n764_));
  XOR2_X1   g563(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n763_), .B(KEYINPUT58), .C1(new_n756_), .C2(new_n757_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n766_), .A2(new_n534_), .A3(new_n538_), .A4(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n762_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n598_), .B1(new_n746_), .B2(new_n752_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(KEYINPUT118), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT118), .B1(new_n770_), .B2(new_n771_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n670_), .B1(new_n769_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n591_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n539_), .A2(new_n571_), .A3(new_n776_), .A4(new_n440_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT54), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n594_), .A2(new_n387_), .A3(new_n608_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G113gat), .B1(new_n782_), .B2(new_n591_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n770_), .A2(new_n771_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n768_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n762_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n784_), .B2(new_n768_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n670_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT122), .B(new_n670_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n778_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n780_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(KEYINPUT123), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT123), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n777_), .B(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n795_), .B1(new_n803_), .B2(new_n792_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n794_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n800_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n799_), .A2(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n591_), .A2(G113gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n783_), .B1(new_n807_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n575_), .B2(KEYINPUT60), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n782_), .B(new_n811_), .C1(KEYINPUT60), .C2(new_n810_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n804_), .A2(new_n575_), .A3(new_n805_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n810_), .ZN(G1341gat));
  AOI21_X1  g613(.A(G127gat), .B1(new_n782_), .B2(new_n440_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n440_), .A2(G127gat), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n807_), .B2(new_n817_), .ZN(G1342gat));
  AOI21_X1  g617(.A(G134gat), .B1(new_n782_), .B2(new_n599_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n637_), .A2(G134gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n807_), .B2(new_n820_), .ZN(G1343gat));
  AND2_X1   g620(.A1(new_n779_), .A2(new_n388_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n594_), .A3(new_n650_), .ZN(new_n823_));
  OR3_X1    g622(.A1(new_n823_), .A2(G141gat), .A3(new_n776_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G141gat), .B1(new_n823_), .B2(new_n776_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1344gat));
  OR3_X1    g625(.A1(new_n823_), .A2(G148gat), .A3(new_n575_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G148gat), .B1(new_n823_), .B2(new_n575_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1345gat));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n823_), .A2(new_n670_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n823_), .B2(new_n670_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1346gat));
  OAI21_X1  g632(.A(G162gat), .B1(new_n823_), .B2(new_n539_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n598_), .A2(G162gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n823_), .B2(new_n835_), .ZN(G1347gat));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n650_), .A2(new_n594_), .A3(new_n663_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n840_), .B2(new_n776_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(KEYINPUT124), .A3(new_n591_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n405_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n793_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n837_), .B1(new_n844_), .B2(G169gat), .ZN(new_n845_));
  AOI211_X1 g644(.A(KEYINPUT62), .B(new_n262_), .C1(new_n793_), .C2(new_n843_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n793_), .A2(new_n626_), .A3(new_n839_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n591_), .A2(new_n273_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT125), .ZN(new_n849_));
  OAI22_X1  g648(.A1(new_n845_), .A2(new_n846_), .B1(new_n847_), .B2(new_n849_), .ZN(G1348gat));
  INV_X1    g649(.A(KEYINPUT126), .ZN(new_n851_));
  INV_X1    g650(.A(new_n271_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n839_), .A2(new_n626_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n803_), .B2(new_n792_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n575_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n852_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n405_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n840_), .A2(new_n263_), .A3(new_n575_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n851_), .B1(new_n856_), .B2(new_n860_), .ZN(new_n861_));
  AOI211_X1 g660(.A(new_n575_), .B(new_n853_), .C1(new_n803_), .C2(new_n792_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT126), .B(new_n859_), .C1(new_n862_), .C2(new_n852_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1349gat));
  NOR3_X1   g663(.A1(new_n847_), .A2(new_n258_), .A3(new_n670_), .ZN(new_n865_));
  INV_X1    g664(.A(G183gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n857_), .A2(new_n440_), .A3(new_n839_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1350gat));
  OAI21_X1  g667(.A(G190gat), .B1(new_n847_), .B2(new_n539_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n854_), .A2(new_n259_), .A3(new_n599_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1351gat));
  NOR2_X1   g670(.A1(new_n650_), .A2(new_n251_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n779_), .A2(new_n388_), .A3(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n776_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n287_), .ZN(G1352gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n575_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n284_), .ZN(G1353gat));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n440_), .B1(new_n879_), .B2(new_n413_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n822_), .A2(new_n878_), .A3(new_n872_), .A4(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT127), .B1(new_n873_), .B2(new_n880_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n413_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n882_), .A2(new_n883_), .A3(new_n879_), .A4(new_n413_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1354gat));
  OAI21_X1  g687(.A(G218gat), .B1(new_n873_), .B2(new_n539_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n598_), .A2(G218gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n873_), .B2(new_n890_), .ZN(G1355gat));
endmodule


