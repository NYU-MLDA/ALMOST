//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n867_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  AND4_X1   g010(.A1(new_n203_), .A2(new_n206_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT8), .B1(new_n207_), .B2(new_n213_), .ZN(new_n214_));
  OR3_X1    g013(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT7), .ZN(new_n216_));
  OR4_X1    g015(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n203_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n207_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n212_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(new_n214_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G57gat), .B(G64gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT11), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(KEYINPUT11), .ZN(new_n224_));
  XOR2_X1   g023(.A(G71gat), .B(G78gat), .Z(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n220_), .A2(new_n221_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT12), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(KEYINPUT12), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G230gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n231_), .A2(new_n232_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n235_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G120gat), .B(G148gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT5), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G176gat), .B(G204gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n240_), .B(new_n241_), .Z(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n238_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT68), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(new_n238_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n242_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT68), .A3(new_n244_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n247_), .A2(new_n249_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT70), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(new_n251_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G1gat), .B(G8gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT73), .ZN(new_n262_));
  INV_X1    g061(.A(G15gat), .ZN(new_n263_));
  INV_X1    g062(.A(G22gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G15gat), .A2(G22gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G1gat), .A2(G8gat), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n265_), .A2(new_n266_), .B1(KEYINPUT14), .B2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n262_), .A2(new_n268_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G29gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G43gat), .B(G50gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n275_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G229gat), .A2(G233gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n275_), .B(KEYINPUT15), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n284_), .A2(new_n271_), .A3(KEYINPUT74), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT74), .B1(new_n284_), .B2(new_n271_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n278_), .A3(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n282_), .B1(new_n287_), .B2(new_n281_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G113gat), .B(G141gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT75), .ZN(new_n290_));
  XOR2_X1   g089(.A(G169gat), .B(G197gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n288_), .B(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n260_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G155gat), .B(G162gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297_));
  INV_X1    g096(.A(G141gat), .ZN(new_n298_));
  INV_X1    g097(.A(G148gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT84), .B1(new_n298_), .B2(new_n299_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G141gat), .A3(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n296_), .B1(new_n304_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n296_), .A2(KEYINPUT1), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n298_), .A2(new_n299_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n305_), .A2(new_n307_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(G228gat), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G78gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(new_n205_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n320_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT87), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(KEYINPUT21), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT21), .ZN(new_n334_));
  INV_X1    g133(.A(new_n331_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n328_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n333_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n317_), .B2(new_n316_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G22gat), .B(G50gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n327_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n327_), .A2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT25), .B(G183gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT24), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n347_), .A2(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G169gat), .ZN(new_n352_));
  INV_X1    g151(.A(G176gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n354_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT76), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n360_), .A3(KEYINPUT23), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362_));
  AND2_X1   g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n358_), .A2(new_n360_), .A3(new_n362_), .A4(KEYINPUT23), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G183gat), .ZN(new_n369_));
  INV_X1    g168(.A(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT23), .B1(new_n358_), .B2(new_n360_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n363_), .A2(new_n364_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G169gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n354_), .B1(new_n375_), .B2(new_n353_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n356_), .A2(new_n368_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT20), .B1(new_n377_), .B2(new_n337_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n366_), .A2(new_n371_), .A3(new_n367_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT78), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G169gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(KEYINPUT78), .A3(new_n352_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n386_));
  AOI21_X1  g185(.A(G176gat), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n354_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n379_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n351_), .B(new_n355_), .C1(new_n373_), .C2(new_n372_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n378_), .B1(new_n394_), .B2(new_n337_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n346_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n377_), .A2(new_n337_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT20), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n338_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT88), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n404_), .B(new_n338_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n399_), .B1(new_n406_), .B2(new_n398_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n389_), .A2(new_n391_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT80), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n404_), .B1(new_n412_), .B2(new_n338_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n405_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n408_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n346_), .A3(new_n397_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G8gat), .B(G36gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n407_), .A2(new_n416_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT96), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n398_), .B(new_n408_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n395_), .A2(new_n398_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n421_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n407_), .A2(new_n416_), .A3(KEYINPUT96), .A4(new_n422_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT27), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n427_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n422_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n428_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n428_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n435_), .B1(new_n440_), .B2(new_n429_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT97), .B1(new_n441_), .B2(new_n436_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n345_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n394_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT82), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447_));
  INV_X1    g246(.A(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(new_n263_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n449_), .B(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT31), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT31), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n446_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n412_), .B(new_n444_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G127gat), .B(G134gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G113gat), .B(G120gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n462_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT83), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n462_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n460_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n457_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n460_), .B(new_n469_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n456_), .A3(new_n454_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT91), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G29gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G57gat), .B(G85gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n477_), .A2(new_n479_), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT4), .ZN(new_n489_));
  INV_X1    g288(.A(new_n465_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n463_), .B1(new_n490_), .B2(new_n467_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(new_n466_), .C1(new_n315_), .C2(new_n310_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n464_), .A2(new_n465_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n311_), .A2(new_n314_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n296_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(new_n303_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n489_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G225gat), .A2(G233gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT4), .B1(new_n470_), .B2(new_n501_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n499_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n316_), .B2(new_n469_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n500_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n488_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(KEYINPUT4), .ZN(new_n508_));
  INV_X1    g307(.A(new_n500_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n502_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(new_n487_), .A3(new_n505_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n507_), .A2(KEYINPUT93), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n488_), .B(new_n514_), .C1(new_n503_), .C2(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT95), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n475_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n436_), .B1(new_n430_), .B2(KEYINPUT27), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n345_), .B1(new_n519_), .B2(new_n517_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n472_), .A2(new_n474_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n522_));
  INV_X1    g321(.A(new_n433_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n421_), .A2(KEYINPUT32), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n516_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n407_), .A2(new_n416_), .A3(KEYINPUT32), .A4(new_n421_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n522_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n434_), .A2(new_n428_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n507_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT33), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT33), .ZN(new_n531_));
  INV_X1    g330(.A(new_n504_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n488_), .B1(new_n532_), .B2(new_n509_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n500_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n531_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n530_), .B1(new_n535_), .B2(new_n529_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n344_), .B1(new_n528_), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n527_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n525_), .A2(new_n522_), .A3(new_n526_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n521_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n443_), .A2(new_n518_), .B1(new_n520_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n220_), .A2(new_n221_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n283_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT34), .ZN(new_n545_));
  OAI221_X1 g344(.A(new_n543_), .B1(KEYINPUT35), .B2(new_n545_), .C1(new_n276_), .C2(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT35), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n551_), .B(KEYINPUT36), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n554_), .B(KEYINPUT71), .Z(new_n560_));
  NOR2_X1   g359(.A1(new_n548_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT37), .B1(new_n553_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n228_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n272_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT16), .ZN(new_n569_));
  XOR2_X1   g368(.A(G183gat), .B(G211gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n566_), .A2(new_n567_), .A3(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(KEYINPUT17), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n566_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n563_), .A2(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n295_), .A2(new_n541_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(G1gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n517_), .B(KEYINPUT98), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT38), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(KEYINPUT100), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(KEYINPUT100), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  NOR2_X1   g383(.A1(new_n295_), .A2(new_n541_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n574_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n557_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n517_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G1gat), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT99), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(new_n591_), .ZN(G1324gat));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n432_), .B1(new_n431_), .B2(new_n437_), .ZN(new_n594_));
  AOI211_X1 g393(.A(KEYINPUT97), .B(new_n436_), .C1(new_n430_), .C2(KEYINPUT27), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n585_), .A2(new_n596_), .A3(new_n587_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(KEYINPUT101), .A3(G8gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT101), .B1(new_n597_), .B2(G8gat), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT102), .B(new_n593_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n600_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n593_), .A2(KEYINPUT102), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n593_), .A2(KEYINPUT102), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n602_), .A2(new_n598_), .A3(new_n603_), .A4(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(G8gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n576_), .A2(new_n606_), .A3(new_n596_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n601_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT40), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n601_), .A2(new_n605_), .A3(KEYINPUT40), .A4(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1325gat));
  OAI21_X1  g411(.A(G15gat), .B1(new_n588_), .B2(new_n475_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT41), .Z(new_n614_));
  NAND3_X1  g413(.A1(new_n576_), .A2(new_n263_), .A3(new_n521_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1326gat));
  OAI21_X1  g415(.A(G22gat), .B1(new_n588_), .B2(new_n344_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT42), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n576_), .A2(new_n264_), .A3(new_n345_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1327gat));
  NOR3_X1   g419(.A1(new_n553_), .A2(new_n556_), .A3(new_n574_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n585_), .A2(new_n621_), .ZN(new_n622_));
  OR3_X1    g421(.A1(new_n622_), .A2(G29gat), .A3(new_n589_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT43), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n344_), .B(new_n518_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n540_), .A2(new_n520_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n563_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AOI211_X1 g428(.A(KEYINPUT43), .B(new_n563_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n294_), .B(new_n586_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT43), .B1(new_n541_), .B2(new_n563_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n627_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n636_), .A2(KEYINPUT44), .A3(new_n294_), .A4(new_n586_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n579_), .A3(new_n637_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n638_), .A2(KEYINPUT103), .A3(G29gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT103), .B1(new_n638_), .B2(G29gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n623_), .B1(new_n639_), .B2(new_n640_), .ZN(G1328gat));
  XOR2_X1   g440(.A(new_n596_), .B(KEYINPUT104), .Z(new_n642_));
  NOR3_X1   g441(.A1(new_n622_), .A2(G36gat), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT45), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n633_), .A2(new_n596_), .A3(new_n637_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G36gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n647_), .A3(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  NOR2_X1   g451(.A1(new_n475_), .A2(new_n448_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n633_), .A2(new_n637_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n633_), .A2(new_n637_), .A3(KEYINPUT105), .A4(new_n653_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n448_), .B1(new_n622_), .B2(new_n475_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .A4(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1330gat));
  AND2_X1   g463(.A1(new_n633_), .A2(new_n637_), .ZN(new_n665_));
  INV_X1    g464(.A(G50gat), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n344_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n585_), .A2(new_n345_), .A3(new_n621_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n665_), .A2(new_n667_), .B1(new_n666_), .B2(new_n668_), .ZN(G1331gat));
  INV_X1    g468(.A(new_n293_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n260_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n541_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n574_), .A3(new_n563_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT107), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(KEYINPUT107), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n579_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(G57gat), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n672_), .A2(new_n587_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n589_), .A2(new_n677_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n676_), .A2(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(G1332gat));
  INV_X1    g479(.A(G64gat), .ZN(new_n681_));
  INV_X1    g480(.A(new_n642_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n678_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n642_), .A2(G64gat), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT109), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n673_), .B2(new_n687_), .ZN(G1333gat));
  INV_X1    g487(.A(G71gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n678_), .B2(new_n521_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT49), .Z(new_n691_));
  NOR2_X1   g490(.A1(new_n475_), .A2(G71gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT110), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n673_), .B2(new_n693_), .ZN(G1334gat));
  AOI21_X1  g493(.A(new_n324_), .B1(new_n678_), .B2(new_n345_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT50), .Z(new_n696_));
  NAND2_X1  g495(.A1(new_n345_), .A2(new_n324_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT111), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n673_), .B2(new_n698_), .ZN(G1335gat));
  NAND2_X1  g498(.A1(new_n672_), .A2(new_n621_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT112), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n209_), .A3(new_n579_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n254_), .A2(new_n259_), .A3(new_n293_), .A4(new_n586_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT114), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(KEYINPUT114), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n636_), .A2(KEYINPUT113), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n636_), .A2(KEYINPUT113), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n517_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n703_), .B1(new_n712_), .B2(new_n209_), .ZN(G1336gat));
  NAND3_X1  g512(.A1(new_n702_), .A2(new_n210_), .A3(new_n596_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n711_), .A2(new_n682_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n210_), .ZN(G1337gat));
  INV_X1    g515(.A(KEYINPUT115), .ZN(new_n717_));
  INV_X1    g516(.A(G99gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n711_), .B2(new_n521_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n521_), .A2(new_n204_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n702_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n717_), .B(KEYINPUT51), .C1(new_n719_), .C2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n717_), .A2(KEYINPUT51), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n475_), .B(new_n708_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n724_), .B(new_n721_), .C1(new_n725_), .C2(new_n718_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1338gat));
  INV_X1    g526(.A(KEYINPUT117), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n704_), .A2(KEYINPUT114), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n344_), .B1(new_n729_), .B2(new_n705_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n205_), .B1(new_n636_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n731_), .A2(KEYINPUT116), .A3(new_n732_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n732_), .A3(G106gat), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n345_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT117), .B(KEYINPUT52), .C1(new_n740_), .C2(new_n205_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n733_), .A2(new_n734_), .A3(new_n738_), .A4(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n702_), .A2(new_n205_), .A3(new_n345_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1339gat));
  INV_X1    g546(.A(G113gat), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n293_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT58), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n237_), .B(KEYINPUT119), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n231_), .A2(new_n232_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n235_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT55), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n754_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n243_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n292_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n280_), .B2(new_n287_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n282_), .B(new_n292_), .C1(new_n287_), .C2(new_n281_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(new_n244_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n750_), .B1(new_n760_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n755_), .A2(new_n756_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n242_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n770_), .A2(KEYINPUT58), .A3(new_n759_), .A4(new_n765_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(new_n628_), .A3(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n758_), .B1(new_n757_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n670_), .A2(new_n244_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n255_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n764_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n557_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n772_), .B1(new_n781_), .B2(KEYINPUT57), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n783_), .B(new_n557_), .C1(new_n778_), .C2(new_n780_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n586_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n575_), .A2(new_n670_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n257_), .A2(new_n251_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n578_), .B1(new_n785_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n443_), .A2(new_n521_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(KEYINPUT59), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT59), .B1(new_n793_), .B2(new_n795_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n749_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n757_), .A2(new_n774_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n776_), .B1(new_n801_), .B2(KEYINPUT56), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n802_), .A2(new_n775_), .B1(new_n779_), .B2(new_n764_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n783_), .B1(new_n803_), .B2(new_n557_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n781_), .A2(KEYINPUT57), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n772_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n791_), .B1(new_n806_), .B2(new_n586_), .ZN(new_n807_));
  NOR4_X1   g606(.A1(new_n807_), .A2(new_n293_), .A3(new_n578_), .A4(new_n794_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n800_), .B1(new_n808_), .B2(G113gat), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n793_), .A2(new_n795_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT121), .B(new_n748_), .C1(new_n810_), .C2(new_n293_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n799_), .A2(new_n809_), .A3(new_n811_), .ZN(G1340gat));
  INV_X1    g611(.A(new_n810_), .ZN(new_n813_));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n671_), .B2(KEYINPUT60), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n813_), .B(new_n815_), .C1(KEYINPUT60), .C2(new_n814_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n798_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n671_), .B1(new_n817_), .B2(new_n796_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n818_), .B2(new_n814_), .ZN(G1341gat));
  INV_X1    g618(.A(G127gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n586_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n822_));
  NOR4_X1   g621(.A1(new_n807_), .A2(new_n586_), .A3(new_n578_), .A4(new_n794_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT122), .B1(new_n823_), .B2(G127gat), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n820_), .C1(new_n810_), .C2(new_n586_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n822_), .A2(new_n824_), .A3(new_n826_), .ZN(G1342gat));
  INV_X1    g626(.A(G134gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n813_), .A2(new_n828_), .A3(new_n557_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n563_), .B1(new_n817_), .B2(new_n796_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n828_), .ZN(G1343gat));
  NOR2_X1   g630(.A1(new_n521_), .A2(new_n344_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n682_), .A2(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n793_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n670_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n260_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g638(.A1(new_n793_), .A2(new_n574_), .A3(new_n834_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT123), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n793_), .A2(new_n842_), .A3(new_n574_), .A4(new_n834_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT61), .B(G155gat), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n841_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1346gat));
  INV_X1    g646(.A(G162gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n835_), .A2(new_n848_), .A3(new_n557_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n835_), .A2(new_n628_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n848_), .ZN(G1347gat));
  XNOR2_X1  g650(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n785_), .A2(new_n792_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n682_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n579_), .A2(new_n345_), .A3(new_n475_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n854_), .A2(new_n293_), .A3(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n852_), .B1(new_n857_), .B2(new_n352_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n852_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n807_), .A2(new_n642_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n855_), .ZN(new_n861_));
  OAI211_X1 g660(.A(G169gat), .B(new_n859_), .C1(new_n861_), .C2(new_n293_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n375_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n858_), .A2(new_n862_), .A3(new_n863_), .ZN(G1348gat));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n260_), .A3(new_n855_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g665(.A1(new_n860_), .A2(new_n574_), .A3(new_n855_), .ZN(new_n867_));
  MUX2_X1   g666(.A(new_n347_), .B(G183gat), .S(new_n867_), .Z(G1350gat));
  AND2_X1   g667(.A1(new_n557_), .A2(new_n348_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n853_), .A2(new_n682_), .A3(new_n855_), .A4(new_n869_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n807_), .A2(new_n563_), .A3(new_n642_), .A4(new_n856_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n370_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT125), .B(new_n870_), .C1(new_n871_), .C2(new_n370_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1351gat));
  NOR2_X1   g675(.A1(new_n833_), .A2(new_n517_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n860_), .A2(new_n670_), .A3(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g678(.A1(new_n854_), .A2(new_n517_), .A3(new_n833_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(G204gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(G204gat), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n880_), .B(new_n260_), .C1(new_n882_), .C2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n860_), .A2(new_n877_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n671_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n886_), .B2(new_n883_), .ZN(G1353gat));
  NAND4_X1  g686(.A1(new_n853_), .A2(new_n574_), .A3(new_n682_), .A4(new_n877_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT63), .B(G211gat), .Z(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  OR3_X1    g689(.A1(new_n888_), .A2(KEYINPUT127), .A3(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n888_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT127), .B1(new_n888_), .B2(new_n890_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n891_), .B1(new_n893_), .B2(new_n894_), .ZN(G1354gat));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n880_), .A2(new_n896_), .A3(new_n557_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G218gat), .B1(new_n885_), .B2(new_n563_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1355gat));
endmodule


