//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(G190gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT23), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT85), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT86), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT87), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT22), .B(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n217_), .B2(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n212_), .B(new_n213_), .C1(new_n216_), .C2(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n210_), .A2(KEYINPUT87), .A3(new_n211_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n207_), .A2(KEYINPUT83), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n223_), .B(new_n204_), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  MUX2_X1   g025(.A(new_n225_), .B(KEYINPUT24), .S(new_n226_), .Z(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT82), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n229_), .B1(new_n203_), .B2(KEYINPUT26), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT26), .B(G190gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n228_), .B(new_n230_), .C1(new_n231_), .C2(new_n229_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  OAI22_X1  g032(.A1(new_n221_), .A2(new_n222_), .B1(new_n224_), .B2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G211gat), .B(G218gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT97), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT96), .B(G204gat), .ZN(new_n237_));
  INV_X1    g036(.A(G197gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G197gat), .A2(G204gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT21), .A3(new_n240_), .ZN(new_n241_));
  MUX2_X1   g040(.A(G204gat), .B(new_n237_), .S(G197gat), .Z(new_n242_));
  OAI211_X1 g041(.A(new_n236_), .B(new_n241_), .C1(KEYINPUT21), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(KEYINPUT21), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n236_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n234_), .A2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT101), .Z(new_n247_));
  XOR2_X1   g046(.A(new_n214_), .B(KEYINPUT99), .Z(new_n248_));
  OAI221_X1 g047(.A(new_n213_), .B1(new_n248_), .B2(G176gat), .C1(new_n211_), .C2(new_n224_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n231_), .A2(new_n228_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n227_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n210_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT20), .B1(new_n252_), .B2(new_n245_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT106), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT19), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n245_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n259_), .B(KEYINPUT20), .C1(new_n234_), .C2(new_n245_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G8gat), .B(G36gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT18), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(KEYINPUT32), .A3(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n253_), .A2(new_n257_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n247_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n260_), .A2(new_n257_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT100), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n260_), .A2(KEYINPUT100), .A3(new_n257_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(KEYINPUT32), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(KEYINPUT104), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT105), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT92), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n282_), .B2(KEYINPUT1), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(KEYINPUT1), .B2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT2), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT93), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(KEYINPUT3), .ZN(new_n291_));
  OR3_X1    g090(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n291_), .B(new_n292_), .C1(new_n288_), .C2(new_n285_), .ZN(new_n293_));
  OAI221_X1 g092(.A(new_n282_), .B1(G155gat), .B2(G162gat), .C1(new_n290_), .C2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT88), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT88), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n296_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n295_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT89), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n304_), .B(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n295_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(new_n312_), .A3(new_n295_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT103), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n308_), .A2(KEYINPUT4), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n314_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n311_), .B1(new_n318_), .B2(new_n310_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G85gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT0), .B(G57gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n266_), .A2(new_n278_), .A3(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n277_), .A2(KEYINPUT105), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT102), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n274_), .A2(new_n331_), .A3(new_n265_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n268_), .A2(new_n265_), .A3(new_n273_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT102), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n332_), .B(new_n334_), .C1(new_n265_), .C2(new_n274_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n325_), .A2(KEYINPUT33), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n318_), .A2(new_n310_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n323_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n336_), .B1(new_n325_), .B2(new_n340_), .ZN(new_n341_));
  OAI22_X1  g140(.A1(new_n329_), .A2(new_n330_), .B1(new_n335_), .B2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n287_), .A2(new_n294_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n345_), .B(KEYINPUT28), .ZN(new_n350_));
  INV_X1    g149(.A(new_n348_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT98), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n349_), .A2(new_n352_), .A3(KEYINPUT98), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n245_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n358_));
  INV_X1    g157(.A(G78gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G106gat), .ZN(new_n361_));
  INV_X1    g160(.A(G228gat), .ZN(new_n362_));
  INV_X1    g161(.A(G233gat), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT94), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(KEYINPUT94), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT95), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n361_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n368_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n357_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G106gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n360_), .B(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n374_), .A2(new_n367_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n369_), .A2(new_n375_), .A3(new_n355_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G43gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n234_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(G15gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT30), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n380_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT91), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n307_), .B(KEYINPUT31), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n387_), .B(KEYINPUT90), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n380_), .A2(new_n384_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n380_), .A2(new_n384_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n387_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(new_n388_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT91), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n377_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n396_), .ZN(new_n399_));
  OAI22_X1  g198(.A1(new_n372_), .A2(new_n376_), .B1(new_n399_), .B2(new_n393_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n355_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n370_), .A2(new_n371_), .A3(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n355_), .B(new_n356_), .C1(new_n369_), .C2(new_n375_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n394_), .A4(new_n396_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n328_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT27), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n333_), .A2(KEYINPUT27), .ZN(new_n407_));
  INV_X1    g206(.A(new_n265_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n261_), .A2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n335_), .A2(new_n406_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n342_), .A2(new_n398_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G229gat), .A2(G233gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G8gat), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(KEYINPUT78), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(KEYINPUT78), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G15gat), .B(G22gat), .ZN(new_n417_));
  INV_X1    g216(.A(G1gat), .ZN(new_n418_));
  INV_X1    g217(.A(G8gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT14), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n414_), .A2(new_n420_), .A3(new_n417_), .A4(new_n415_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G29gat), .B(G36gat), .Z(new_n425_));
  XOR2_X1   g224(.A(G43gat), .B(G50gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n422_), .A2(new_n423_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n427_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n412_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n427_), .B(KEYINPUT15), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n424_), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n412_), .B(KEYINPUT81), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(new_n430_), .B2(new_n427_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n432_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G113gat), .B(G141gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G169gat), .B(G197gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n438_), .B(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G230gat), .A2(G233gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT65), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT66), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT65), .B1(KEYINPUT66), .B2(KEYINPUT7), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G99gat), .A2(G106gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT64), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n458_), .A2(KEYINPUT64), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n455_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n455_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(KEYINPUT64), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n450_), .A2(new_n454_), .B1(new_n460_), .B2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G85gat), .B(G92gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT8), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n464_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT7), .B1(new_n447_), .B2(KEYINPUT66), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n373_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n451_), .ZN(new_n474_));
  OAI22_X1  g273(.A1(new_n469_), .A2(new_n470_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT8), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n466_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n468_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G71gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(G78gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n359_), .A2(G71gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G57gat), .B(G64gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(KEYINPUT11), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT67), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n483_), .B2(KEYINPUT11), .ZN(new_n486_));
  INV_X1    g285(.A(G64gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G57gat), .ZN(new_n488_));
  INV_X1    g287(.A(G57gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G64gat), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n488_), .A2(new_n490_), .A3(new_n485_), .A4(KEYINPUT11), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n484_), .B1(new_n486_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n488_), .A2(new_n490_), .A3(KEYINPUT11), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT67), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n490_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n495_), .A2(new_n498_), .A3(new_n482_), .A4(new_n491_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n493_), .A2(new_n499_), .A3(KEYINPUT68), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n499_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT68), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G85gat), .ZN(new_n504_));
  INV_X1    g303(.A(G92gat), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT9), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n466_), .B2(KEYINPUT9), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n460_), .A2(new_n464_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT10), .B(G99gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(G106gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n478_), .A2(new_n500_), .A3(new_n503_), .A4(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n493_), .A2(new_n499_), .A3(KEYINPUT68), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT68), .B1(new_n493_), .B2(new_n499_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n511_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n468_), .B2(new_n477_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n445_), .B1(new_n513_), .B2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n473_), .B2(new_n446_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n454_), .B1(new_n524_), .B2(KEYINPUT7), .ZN(new_n525_));
  AOI211_X1 g324(.A(KEYINPUT8), .B(new_n467_), .C1(new_n525_), .C2(new_n508_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n476_), .B1(new_n475_), .B2(new_n466_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n511_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n493_), .A2(new_n499_), .A3(KEYINPUT12), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n522_), .A2(new_n444_), .A3(new_n512_), .A4(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G120gat), .B(G148gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT70), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n532_), .B(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n539_), .A2(KEYINPUT13), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(KEYINPUT13), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT75), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT34), .Z(new_n546_));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n546_), .A2(new_n547_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT74), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n551_), .B1(new_n528_), .B2(new_n433_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n528_), .A2(KEYINPUT72), .A3(new_n428_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n518_), .B2(new_n427_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n552_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n550_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT72), .B1(new_n528_), .B2(new_n428_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n518_), .A2(new_n554_), .A3(new_n427_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n557_), .B1(new_n562_), .B2(new_n552_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT73), .ZN(new_n566_));
  XOR2_X1   g365(.A(G134gat), .B(G162gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n544_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n556_), .A2(new_n558_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n562_), .A2(new_n557_), .A3(new_n552_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(KEYINPUT75), .A3(new_n569_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n568_), .B(KEYINPUT36), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n564_), .A2(KEYINPUT76), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n571_), .A2(new_n575_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT77), .B(KEYINPUT37), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT75), .B1(new_n574_), .B2(new_n569_), .ZN(new_n583_));
  AOI211_X1 g382(.A(new_n544_), .B(new_n570_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n584_));
  OAI22_X1  g383(.A1(new_n583_), .A2(new_n584_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT37), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n424_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n503_), .A2(new_n500_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT80), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT17), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n501_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n589_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n600_), .B2(new_n589_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(KEYINPUT17), .B2(new_n597_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n587_), .A2(new_n604_), .ZN(new_n605_));
  NOR4_X1   g404(.A1(new_n411_), .A2(new_n443_), .A3(new_n543_), .A4(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n418_), .A3(new_n328_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n411_), .A2(new_n580_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n604_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n611_), .A2(new_n543_), .A3(new_n443_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n418_), .B1(new_n613_), .B2(new_n328_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n615_), .B1(new_n608_), .B2(new_n607_), .ZN(G1324gat));
  INV_X1    g415(.A(new_n410_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n606_), .A2(new_n419_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G8gat), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(KEYINPUT39), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(KEYINPUT39), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n618_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1325gat));
  AOI21_X1  g424(.A(new_n382_), .B1(new_n613_), .B2(new_n397_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT41), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n606_), .A2(new_n382_), .A3(new_n397_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1326gat));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n613_), .B2(new_n377_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT42), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n377_), .A2(new_n630_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT107), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n606_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(G1327gat));
  NOR2_X1   g435(.A1(new_n411_), .A2(new_n443_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n611_), .A2(new_n580_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n543_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n328_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT43), .B1(new_n411_), .B2(new_n587_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n342_), .A2(new_n398_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n405_), .A2(new_n410_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n580_), .A2(new_n581_), .B1(new_n585_), .B2(KEYINPUT37), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n643_), .A2(new_n649_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n543_), .A2(new_n443_), .A3(new_n604_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT109), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT108), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n651_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n643_), .B2(new_n649_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n653_), .B1(new_n658_), .B2(KEYINPUT108), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n659_), .B2(KEYINPUT44), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n328_), .A2(G29gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n642_), .B1(new_n660_), .B2(new_n661_), .ZN(G1328gat));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n660_), .B2(new_n617_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n641_), .A2(new_n663_), .A3(new_n617_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT45), .Z(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(new_n668_), .A3(KEYINPUT46), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1329gat));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n650_), .A2(KEYINPUT108), .A3(new_n651_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT44), .B1(new_n674_), .B2(KEYINPUT109), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n652_), .A2(new_n655_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n397_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G43gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n397_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n640_), .A2(G43gat), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n673_), .B1(new_n678_), .B2(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT47), .B(new_n680_), .C1(new_n677_), .C2(G43gat), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1330gat));
  INV_X1    g483(.A(G50gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n641_), .A2(new_n685_), .A3(new_n377_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n660_), .A2(new_n377_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(KEYINPUT110), .ZN(new_n688_));
  OAI21_X1  g487(.A(G50gat), .B1(new_n687_), .B2(KEYINPUT110), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(G1331gat));
  AND4_X1   g489(.A1(new_n443_), .A2(new_n610_), .A3(new_n543_), .A4(new_n604_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(G57gat), .A3(new_n328_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT112), .ZN(new_n693_));
  NOR4_X1   g492(.A1(new_n411_), .A2(new_n442_), .A3(new_n542_), .A4(new_n605_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n328_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT111), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT111), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n693_), .A2(new_n696_), .A3(new_n697_), .ZN(G1332gat));
  AOI21_X1  g497(.A(new_n487_), .B1(new_n691_), .B2(new_n617_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT48), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n694_), .A2(new_n487_), .A3(new_n617_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1333gat));
  AOI21_X1  g501(.A(new_n479_), .B1(new_n691_), .B2(new_n397_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n694_), .A2(new_n479_), .A3(new_n397_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1334gat));
  AOI21_X1  g506(.A(new_n359_), .B1(new_n691_), .B2(new_n377_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT50), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n694_), .A2(new_n359_), .A3(new_n377_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1335gat));
  NAND3_X1  g510(.A1(new_n611_), .A2(new_n543_), .A3(new_n443_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT114), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n643_), .B2(new_n649_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n328_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G85gat), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NOR4_X1   g516(.A1(new_n411_), .A2(new_n442_), .A3(new_n542_), .A4(new_n638_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n504_), .A3(new_n328_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1336gat));
  OAI21_X1  g519(.A(G92gat), .B1(new_n715_), .B2(new_n410_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n505_), .A3(new_n617_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1337gat));
  OAI21_X1  g522(.A(G99gat), .B1(new_n715_), .B2(new_n679_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n679_), .A2(new_n509_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n718_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g527(.A1(new_n718_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n714_), .A2(new_n377_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G106gat), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT52), .B(new_n373_), .C1(new_n714_), .C2(new_n377_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g534(.A1(new_n617_), .A2(new_n716_), .A3(new_n400_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n539_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n434_), .A2(new_n431_), .A3(new_n436_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n429_), .A2(new_n431_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n441_), .B1(new_n740_), .B2(new_n435_), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n438_), .A2(new_n441_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n530_), .A2(new_n512_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n521_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n590_), .B2(new_n528_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n522_), .A2(KEYINPUT115), .A3(new_n512_), .A4(new_n530_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n445_), .A3(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n745_), .A2(new_n747_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(KEYINPUT55), .A4(new_n444_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT116), .B1(new_n531_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n531_), .A2(new_n754_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n750_), .A2(new_n753_), .A3(new_n755_), .A4(new_n756_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n537_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(KEYINPUT117), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n537_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(KEYINPUT117), .A3(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n532_), .A2(new_n537_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n442_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n743_), .B1(new_n760_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n580_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(KEYINPUT57), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  INV_X1    g570(.A(new_n743_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n761_), .A2(new_n762_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n765_), .B1(new_n759_), .B2(KEYINPUT117), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n772_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n771_), .B1(new_n778_), .B2(new_n580_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n764_), .A2(new_n742_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT58), .B(new_n780_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n773_), .A2(new_n775_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(KEYINPUT118), .A3(KEYINPUT58), .A4(new_n780_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n780_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n783_), .A2(new_n785_), .A3(new_n788_), .A4(new_n648_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n770_), .A2(new_n779_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n611_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n587_), .A2(new_n443_), .A3(new_n542_), .A4(new_n604_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT54), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT119), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(new_n793_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n737_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(G113gat), .B1(new_n798_), .B2(new_n442_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n797_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n796_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n736_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n737_), .A2(KEYINPUT59), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n802_), .A2(new_n806_), .B1(new_n794_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(G113gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n442_), .B2(KEYINPUT121), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(KEYINPUT121), .B2(new_n809_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n799_), .B1(new_n808_), .B2(new_n811_), .ZN(G1340gat));
  INV_X1    g611(.A(G120gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n542_), .B2(KEYINPUT60), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n798_), .B(new_n814_), .C1(KEYINPUT60), .C2(new_n813_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n794_), .A2(new_n736_), .A3(new_n801_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n543_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n802_), .B2(new_n806_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G120gat), .B1(new_n818_), .B2(KEYINPUT122), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT122), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n817_), .C1(new_n802_), .C2(new_n806_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT123), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n815_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n808_), .B2(new_n604_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n798_), .A2(new_n827_), .A3(new_n604_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n828_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n808_), .A2(new_n648_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G134gat), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n769_), .A2(G134gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n805_), .B2(new_n837_), .ZN(G1343gat));
  AOI21_X1  g637(.A(new_n404_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n410_), .A3(new_n328_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n443_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT125), .B(G141gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1344gat));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n542_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT126), .B(G148gat), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1345gat));
  NOR2_X1   g645(.A1(new_n840_), .A2(new_n611_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT61), .B(G155gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  OAI21_X1  g648(.A(G162gat), .B1(new_n840_), .B2(new_n587_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n769_), .A2(G162gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n840_), .B2(new_n851_), .ZN(G1347gat));
  NOR3_X1   g651(.A1(new_n410_), .A2(new_n328_), .A3(new_n400_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n794_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n442_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n855_), .B(G169gat), .C1(KEYINPUT127), .C2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT127), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(KEYINPUT62), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(KEYINPUT127), .A3(new_n856_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n860_), .B(new_n861_), .C1(new_n248_), .C2(new_n855_), .ZN(G1348gat));
  AOI21_X1  g661(.A(G176gat), .B1(new_n854_), .B2(new_n543_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n377_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n410_), .A2(new_n328_), .ZN(new_n865_));
  AND4_X1   g664(.A1(G176gat), .A2(new_n865_), .A3(new_n397_), .A4(new_n543_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n864_), .B2(new_n866_), .ZN(G1349gat));
  INV_X1    g666(.A(new_n854_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(new_n228_), .A3(new_n611_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n864_), .A2(new_n397_), .A3(new_n604_), .A4(new_n865_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n202_), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n868_), .B2(new_n587_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n854_), .A2(new_n231_), .A3(new_n580_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1351gat));
  NAND2_X1  g673(.A1(new_n839_), .A2(new_n865_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n443_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n238_), .ZN(G1352gat));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n542_), .ZN(new_n878_));
  MUX2_X1   g677(.A(G204gat), .B(new_n237_), .S(new_n878_), .Z(G1353gat));
  NOR2_X1   g678(.A1(new_n875_), .A2(new_n611_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n880_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT63), .B(G211gat), .Z(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n880_), .B2(new_n882_), .ZN(G1354gat));
  OAI21_X1  g682(.A(G218gat), .B1(new_n875_), .B2(new_n587_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n769_), .A2(G218gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n875_), .B2(new_n885_), .ZN(G1355gat));
endmodule


