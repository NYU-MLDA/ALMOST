//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n211_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  MUX2_X1   g013(.A(new_n204_), .B(new_n205_), .S(new_n214_), .Z(new_n215_));
  NAND2_X1  g014(.A1(G229gat), .A2(G233gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n215_), .A2(KEYINPUT78), .A3(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n214_), .B(new_n204_), .Z(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT78), .B1(new_n215_), .B2(new_n217_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G141gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G169gat), .B(G197gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n227_), .B(KEYINPUT79), .Z(new_n228_));
  OR2_X1    g027(.A1(new_n222_), .A2(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT6), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  OR3_X1    g033(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT8), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n236_), .A2(new_n241_), .A3(new_n237_), .A4(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT10), .B(G99gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT64), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT65), .B(G106gat), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n238_), .A2(KEYINPUT9), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT67), .B(G92gat), .ZN(new_n250_));
  INV_X1    g049(.A(G85gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT9), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n249_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n237_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n233_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n246_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n243_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT68), .B(G71gat), .ZN(new_n258_));
  INV_X1    g057(.A(G78gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G57gat), .B(G64gat), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(KEYINPUT11), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(KEYINPUT11), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n260_), .B1(new_n264_), .B2(new_n262_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n257_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n257_), .A2(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G230gat), .A2(G233gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n257_), .A2(KEYINPUT69), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n243_), .B(new_n274_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n273_), .A2(KEYINPUT12), .A3(new_n275_), .A4(new_n266_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n267_), .A2(new_n270_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(G230gat), .A3(G233gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G120gat), .B(G148gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT5), .ZN(new_n282_));
  XOR2_X1   g081(.A(G176gat), .B(G204gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(KEYINPUT71), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(KEYINPUT13), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(KEYINPUT13), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n231_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  OR2_X1    g093(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n295_), .A2(KEYINPUT89), .A3(G197gat), .A4(new_n296_), .ZN(new_n297_));
  AND2_X1   g096(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n299_));
  INV_X1    g098(.A(G197gat), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G204gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT89), .B1(new_n302_), .B2(G197gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n294_), .B(new_n297_), .C1(new_n301_), .C2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT90), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT88), .B(G204gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n303_), .B1(new_n308_), .B2(new_n300_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n309_), .A2(KEYINPUT90), .A3(new_n294_), .A4(new_n297_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G211gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(G218gat), .ZN(new_n313_));
  INV_X1    g112(.A(G218gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n314_), .A2(G211gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n300_), .A2(G204gat), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n308_), .B2(new_n300_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n318_), .B2(new_n294_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n311_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT85), .A4(new_n326_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n329_), .A2(new_n330_), .B1(G169gat), .B2(G176gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n332_));
  NAND2_X1  g131(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n332_), .B(G169gat), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT84), .B(G176gat), .ZN(new_n337_));
  INV_X1    g136(.A(G169gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n335_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n333_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT83), .B1(new_n338_), .B2(KEYINPUT22), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n336_), .B(new_n337_), .C1(new_n340_), .C2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT24), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT25), .B(G183gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT80), .B1(new_n348_), .B2(G190gat), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT26), .B(G190gat), .Z(new_n351_));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n346_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT24), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n345_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT81), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n356_), .A2(new_n324_), .A3(KEYINPUT81), .A4(new_n326_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n331_), .A2(new_n342_), .B1(new_n354_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n297_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT21), .B1(new_n313_), .B2(new_n315_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT91), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT91), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n321_), .A2(new_n362_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n337_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT22), .B(G169gat), .Z(new_n373_));
  OAI211_X1 g172(.A(new_n327_), .B(new_n343_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT26), .B(G190gat), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n375_), .A2(new_n347_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n376_), .A2(new_n357_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n344_), .B(KEYINPUT96), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(new_n345_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n374_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  AOI211_X1 g179(.A(KEYINPUT91), .B(new_n364_), .C1(new_n309_), .C2(new_n297_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n368_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n319_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n380_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n371_), .A2(new_n385_), .A3(KEYINPUT20), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT18), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n321_), .A2(new_n380_), .A3(new_n370_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n362_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n389_), .ZN(new_n399_));
  AND4_X1   g198(.A1(KEYINPUT97), .A2(new_n398_), .A3(KEYINPUT20), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT97), .B1(new_n402_), .B2(new_n399_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n390_), .B(new_n395_), .C1(new_n400_), .C2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n386_), .A2(new_n399_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(KEYINPUT20), .A3(new_n389_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT99), .A4(new_n394_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n394_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT99), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT27), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n390_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n394_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT27), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n404_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G141gat), .A2(G148gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT3), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G141gat), .A2(G148gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT2), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(KEYINPUT1), .B2(new_n423_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(KEYINPUT1), .B2(new_n423_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n418_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n430_), .A2(new_n420_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G127gat), .B(G134gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G113gat), .B(G120gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n433_), .A2(new_n434_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n427_), .B(new_n432_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n427_), .A2(new_n432_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(KEYINPUT87), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n438_), .B(KEYINPUT4), .C1(new_n439_), .C2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n427_), .A2(new_n432_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n444_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n447_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(new_n438_), .A3(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT0), .ZN(new_n456_));
  INV_X1    g255(.A(G57gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(new_n251_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n458_), .B(G85gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n451_), .A2(new_n461_), .A3(new_n453_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n321_), .A2(new_n370_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n447_), .A2(KEYINPUT29), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G228gat), .ZN(new_n467_));
  INV_X1    g266(.A(G233gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT92), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n467_), .A2(new_n468_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n466_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n464_), .A2(new_n471_), .A3(new_n465_), .A4(new_n470_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n447_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT28), .B1(new_n447_), .B2(KEYINPUT29), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G22gat), .B(G50gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n473_), .A2(new_n475_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n476_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT94), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n489_), .A3(new_n486_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT93), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n484_), .A2(new_n488_), .A3(new_n490_), .A4(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n487_), .A2(new_n491_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n463_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n417_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT100), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n417_), .A2(KEYINPUT100), .A3(new_n496_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n395_), .A2(KEYINPUT32), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n413_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n405_), .A2(new_n406_), .A3(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n463_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT98), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT98), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n506_), .B(new_n507_), .C1(new_n413_), .C2(new_n501_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n444_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n452_), .A2(new_n438_), .A3(new_n450_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n459_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT33), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n462_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n512_), .B2(new_n462_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n414_), .A2(new_n514_), .A3(new_n404_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n505_), .A2(new_n508_), .A3(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n493_), .A2(new_n495_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n499_), .A2(new_n500_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n362_), .B(KEYINPUT30), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G71gat), .B(G99gat), .ZN(new_n521_));
  INV_X1    g320(.A(G43gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G227gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(G15gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n523_), .B(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n520_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n362_), .A2(KEYINPUT30), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n362_), .A2(KEYINPUT30), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n527_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT86), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n520_), .A2(new_n533_), .A3(new_n527_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n528_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI211_X1 g336(.A(KEYINPUT31), .B(new_n528_), .C1(new_n532_), .C2(new_n534_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n443_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n532_), .A2(new_n534_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT31), .B1(new_n540_), .B2(new_n528_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n536_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(new_n445_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n463_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n517_), .A2(new_n544_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT101), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n417_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n412_), .A2(KEYINPUT101), .A3(new_n416_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n519_), .A2(new_n545_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n293_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT37), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n273_), .A2(new_n275_), .A3(new_n205_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT74), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT74), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n273_), .A2(new_n557_), .A3(new_n275_), .A4(new_n205_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n257_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n560_), .A2(new_n204_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n559_), .B(new_n565_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(KEYINPUT75), .A3(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G190gat), .B(G218gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n569_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n573_), .A2(new_n574_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n570_), .A2(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n568_), .A2(KEYINPUT75), .A3(new_n569_), .A4(new_n575_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n554_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n570_), .A2(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n578_), .ZN(new_n583_));
  AND4_X1   g382(.A1(new_n554_), .A2(new_n582_), .A3(new_n580_), .A4(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n266_), .B(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n214_), .B(KEYINPUT76), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G127gat), .B(G155gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT16), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT17), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n589_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n589_), .A2(new_n595_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT77), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n585_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n553_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT102), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n463_), .B(KEYINPUT103), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n207_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT105), .Z(new_n609_));
  AND2_X1   g408(.A1(new_n579_), .A2(new_n580_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT104), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT104), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n552_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n599_), .A3(new_n292_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n546_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n609_), .B(new_n616_), .C1(new_n607_), .C2(new_n606_), .ZN(G1324gat));
  INV_X1    g416(.A(new_n550_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT101), .B1(new_n412_), .B2(new_n416_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n603_), .A2(new_n208_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G8gat), .B1(new_n615_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT39), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(G1325gat));
  OAI21_X1  g426(.A(G15gat), .B1(new_n615_), .B2(new_n545_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(KEYINPUT41), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n544_), .A2(new_n525_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n629_), .B(new_n630_), .C1(new_n602_), .C2(new_n631_), .ZN(G1326gat));
  OAI21_X1  g431(.A(G22gat), .B1(new_n615_), .B2(new_n517_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT42), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n517_), .A2(G22gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n602_), .B2(new_n635_), .ZN(G1327gat));
  INV_X1    g435(.A(new_n613_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n600_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n553_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n463_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n581_), .A2(new_n584_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n643_), .B(KEYINPUT43), .C1(new_n552_), .C2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n519_), .A2(new_n545_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n547_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n647_), .B(new_n546_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n644_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT107), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT108), .B1(new_n649_), .B2(new_n650_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT108), .ZN(new_n653_));
  NOR4_X1   g452(.A1(new_n552_), .A2(new_n653_), .A3(KEYINPUT43), .A4(new_n644_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n645_), .B(new_n651_), .C1(new_n652_), .C2(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n655_), .A2(new_n600_), .A3(new_n292_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT44), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(G29gat), .A3(new_n605_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n656_), .A2(KEYINPUT44), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n642_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n657_), .A3(new_n620_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n640_), .A2(G36gat), .A3(new_n622_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT45), .Z(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(KEYINPUT46), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  NAND4_X1  g468(.A1(new_n659_), .A2(new_n657_), .A3(G43gat), .A4(new_n544_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n522_), .B1(new_n640_), .B2(new_n545_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g472(.A1(new_n493_), .A2(new_n495_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G50gat), .B1(new_n641_), .B2(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n657_), .A2(G50gat), .A3(new_n674_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(new_n659_), .ZN(G1331gat));
  INV_X1    g476(.A(new_n552_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n291_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n230_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n601_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n605_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n614_), .A2(new_n638_), .A3(new_n680_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT109), .Z(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT110), .B(G57gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n546_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n685_), .B1(new_n687_), .B2(new_n689_), .ZN(G1332gat));
  INV_X1    g489(.A(G64gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n687_), .B2(new_n620_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT48), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n691_), .A3(new_n620_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1333gat));
  INV_X1    g494(.A(G71gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n687_), .B2(new_n544_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n684_), .A2(new_n696_), .A3(new_n544_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  AOI21_X1  g500(.A(new_n259_), .B1(new_n687_), .B2(new_n674_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n674_), .A2(new_n259_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT113), .Z(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n683_), .B2(new_n706_), .ZN(G1335gat));
  NOR3_X1   g506(.A1(new_n681_), .A2(new_n638_), .A3(new_n637_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n251_), .A3(new_n605_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n680_), .A2(new_n600_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n655_), .A2(KEYINPUT114), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n655_), .A2(KEYINPUT114), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(new_n463_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n714_), .B2(new_n251_), .ZN(G1336gat));
  AOI21_X1  g514(.A(G92gat), .B1(new_n708_), .B2(new_n620_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n622_), .A2(new_n250_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n713_), .B2(new_n717_), .ZN(G1337gat));
  AND3_X1   g517(.A1(new_n708_), .A2(new_n245_), .A3(new_n544_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n544_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(G99gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g521(.A(KEYINPUT115), .ZN(new_n723_));
  INV_X1    g522(.A(new_n645_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n497_), .A2(new_n498_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n544_), .B1(new_n725_), .B2(new_n500_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n648_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n585_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n643_), .B1(new_n728_), .B2(KEYINPUT43), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n724_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n585_), .B(new_n650_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n653_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n649_), .A2(KEYINPUT108), .A3(new_n650_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n638_), .B1(new_n730_), .B2(new_n734_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n230_), .A2(new_n679_), .A3(new_n517_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n723_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n655_), .A2(new_n723_), .A3(new_n600_), .A4(new_n736_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G106gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT52), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT117), .ZN(new_n741_));
  INV_X1    g540(.A(new_n739_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n655_), .A2(new_n600_), .A3(new_n736_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT115), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .A4(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n746_), .A2(new_n744_), .A3(G106gat), .A4(new_n738_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT116), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(KEYINPUT52), .C1(new_n737_), .C2(new_n739_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n741_), .A2(new_n747_), .A3(new_n749_), .A4(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n708_), .A2(new_n247_), .A3(new_n674_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n756_), .A3(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  NAND2_X1  g557(.A1(new_n551_), .A2(new_n605_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT57), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n231_), .A2(new_n285_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n272_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n277_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n277_), .A2(new_n764_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n286_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n762_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n226_), .B1(new_n219_), .B2(new_n216_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n215_), .B(KEYINPUT120), .Z(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n216_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n228_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n288_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n761_), .B(new_n637_), .C1(new_n776_), .C2(new_n782_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n762_), .A2(new_n775_), .B1(new_n781_), .B2(new_n780_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT57), .B1(new_n784_), .B2(new_n613_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n285_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n775_), .A2(new_n787_), .A3(new_n780_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n788_), .A2(KEYINPUT58), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n644_), .B1(new_n788_), .B2(KEYINPUT58), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n599_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n601_), .A2(new_n231_), .A3(new_n679_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n793_), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT118), .B1(new_n793_), .B2(KEYINPUT54), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(KEYINPUT54), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n760_), .B1(new_n792_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(G113gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(new_n230_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n797_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n783_), .A2(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n638_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n759_), .B(KEYINPUT121), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n803_), .A2(new_n810_), .A3(new_n231_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n801_), .B1(new_n811_), .B2(new_n800_), .ZN(G1340gat));
  NAND3_X1  g611(.A1(new_n802_), .A2(new_n291_), .A3(new_n809_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n802_), .A2(KEYINPUT123), .A3(new_n291_), .A4(new_n809_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(G120gat), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n818_));
  AOI21_X1  g617(.A(G120gat), .B1(new_n291_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT122), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n819_), .A2(new_n820_), .B1(new_n818_), .B2(G120gat), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n799_), .B(new_n821_), .C1(new_n820_), .C2(new_n819_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n822_), .ZN(G1341gat));
  INV_X1    g622(.A(G127gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n799_), .A2(new_n824_), .A3(new_n638_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n599_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n803_), .A2(new_n810_), .A3(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n827_), .B2(new_n824_), .ZN(G1342gat));
  INV_X1    g627(.A(G134gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n799_), .A2(new_n829_), .A3(new_n613_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n803_), .A2(new_n810_), .A3(new_n644_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n829_), .ZN(G1343gat));
  INV_X1    g631(.A(new_n792_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n804_), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n620_), .A2(new_n544_), .A3(new_n517_), .A4(new_n604_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n230_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n291_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g640(.A1(new_n836_), .A2(new_n600_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT61), .B(G155gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  OAI21_X1  g643(.A(G162gat), .B1(new_n836_), .B2(new_n644_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n637_), .A2(G162gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n836_), .B2(new_n846_), .ZN(G1347gat));
  NAND3_X1  g646(.A1(new_n620_), .A2(new_n544_), .A3(new_n604_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT124), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n674_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n638_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n230_), .B(new_n850_), .C1(new_n851_), .C2(new_n797_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n373_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n806_), .A2(KEYINPUT125), .A3(new_n230_), .A4(new_n850_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n338_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n853_), .B1(new_n857_), .B2(KEYINPUT62), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(KEYINPUT62), .B2(new_n857_), .ZN(G1348gat));
  AND2_X1   g658(.A1(new_n806_), .A2(new_n850_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n372_), .B1(new_n860_), .B2(new_n291_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n674_), .B1(new_n833_), .B2(new_n804_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n849_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n863_), .A2(G176gat), .A3(new_n291_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n862_), .B2(new_n864_), .ZN(G1349gat));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n638_), .A3(new_n863_), .ZN(new_n866_));
  INV_X1    g665(.A(G183gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n826_), .A2(new_n347_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n866_), .A2(new_n867_), .B1(new_n860_), .B2(new_n868_), .ZN(G1350gat));
  NAND2_X1  g668(.A1(new_n860_), .A2(new_n585_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G190gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n860_), .A2(new_n375_), .A3(new_n613_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1351gat));
  NAND2_X1  g672(.A1(new_n545_), .A2(new_n496_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n620_), .B1(KEYINPUT126), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(KEYINPUT126), .B2(new_n874_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n834_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n231_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n300_), .ZN(G1352gat));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n877_), .A2(new_n679_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n302_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT127), .B(G204gat), .C1(new_n877_), .C2(new_n679_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .ZN(G1353gat));
  INV_X1    g684(.A(new_n877_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT63), .B(G211gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n599_), .A3(new_n887_), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n877_), .A2(new_n826_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1354gat));
  OAI21_X1  g689(.A(G218gat), .B1(new_n877_), .B2(new_n644_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n613_), .A2(new_n314_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n877_), .B2(new_n892_), .ZN(G1355gat));
endmodule


