//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n851_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT37), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT35), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G29gat), .B(G36gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209_));
  OR3_X1    g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n209_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G85gat), .A3(G92gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT9), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(new_n224_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(G99gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n222_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n233_), .A2(new_n215_), .A3(new_n218_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n227_), .A2(new_n228_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n230_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n212_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT15), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n212_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n224_), .A2(new_n229_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(new_n219_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n220_), .A2(KEYINPUT67), .A3(new_n224_), .A4(new_n229_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n235_), .A2(new_n237_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT8), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT66), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n241_), .B1(new_n243_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT34), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(KEYINPUT69), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n256_), .B2(KEYINPUT69), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n204_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n256_), .A2(new_n204_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n260_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G190gat), .B(G218gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(G134gat), .B(G162gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT36), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(new_n266_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n269_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT36), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n203_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n264_), .A2(new_n265_), .A3(new_n260_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT35), .B1(new_n264_), .B2(new_n260_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n274_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n202_), .A2(KEYINPUT37), .ZN(new_n281_));
  INV_X1    g080(.A(new_n203_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n280_), .A2(new_n271_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285_));
  INV_X1    g084(.A(G1gat), .ZN(new_n286_));
  INV_X1    g085(.A(G8gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT14), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G1gat), .B(G8gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G231gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G57gat), .B(G64gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G71gat), .B(G78gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT11), .ZN(new_n296_));
  XOR2_X1   g095(.A(G71gat), .B(G78gat), .Z(new_n297_));
  INV_X1    g096(.A(G64gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G57gat), .ZN(new_n299_));
  INV_X1    g098(.A(G57gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G64gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n301_), .A3(KEYINPUT11), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n294_), .A2(KEYINPUT11), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n296_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n293_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G127gat), .B(G155gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT16), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G183gat), .B(G211gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT17), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(KEYINPUT17), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT71), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n307_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT72), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(KEYINPUT72), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n313_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n284_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT73), .ZN(new_n321_));
  INV_X1    g120(.A(G183gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT77), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT25), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n322_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT78), .ZN(new_n328_));
  XOR2_X1   g127(.A(KEYINPUT26), .B(G190gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(G183gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(KEYINPUT25), .B2(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT23), .ZN(new_n334_));
  OR2_X1    g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT24), .A3(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n334_), .B(new_n337_), .C1(KEYINPUT24), .C2(new_n335_), .ZN(new_n338_));
  INV_X1    g137(.A(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n330_), .A2(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n340_), .A2(new_n334_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n336_), .B1(new_n343_), .B2(G176gat), .ZN(new_n344_));
  OAI22_X1  g143(.A1(new_n332_), .A2(new_n338_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G71gat), .B(G99gat), .ZN(new_n348_));
  INV_X1    g147(.A(G43gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351_));
  INV_X1    g150(.A(G15gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n350_), .B(new_n353_), .Z(new_n354_));
  NAND2_X1  g153(.A1(new_n345_), .A2(new_n346_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n347_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n347_), .B2(new_n355_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT31), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G127gat), .B(G134gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT79), .ZN(new_n361_));
  XOR2_X1   g160(.A(G113gat), .B(G120gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n345_), .B(new_n346_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n354_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n356_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n359_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n359_), .B2(new_n368_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G197gat), .B(G204gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT85), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT21), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT84), .Z(new_n378_));
  NOR2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT21), .ZN(new_n380_));
  INV_X1    g179(.A(G197gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G204gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(new_n373_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n385_), .A2(new_n377_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n379_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G228gat), .ZN(new_n388_));
  INV_X1    g187(.A(G233gat), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G141gat), .ZN(new_n396_));
  INV_X1    g195(.A(G148gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT81), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT2), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n400_), .A2(new_n401_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n396_), .A2(new_n397_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n404_), .B2(new_n402_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n395_), .B1(new_n399_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n392_), .B1(new_n394_), .B2(KEYINPUT1), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(KEYINPUT1), .B2(new_n392_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n396_), .A2(new_n397_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n411_), .A3(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT29), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n387_), .A2(new_n391_), .A3(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n379_), .A2(new_n386_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT86), .B1(new_n379_), .B2(new_n386_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n418_), .A2(new_n419_), .B1(KEYINPUT29), .B2(new_n413_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n415_), .B1(new_n420_), .B2(new_n391_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n415_), .B(new_n424_), .C1(new_n420_), .C2(new_n391_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n426_));
  AND3_X1   g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n413_), .A2(KEYINPUT29), .ZN(new_n429_));
  XOR2_X1   g228(.A(G22gat), .B(G50gat), .Z(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n427_), .A2(new_n428_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n418_), .A2(new_n419_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n414_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n390_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n424_), .B1(new_n437_), .B2(new_n415_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n425_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n434_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n431_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n372_), .B1(new_n433_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n359_), .A2(new_n368_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n363_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n369_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n432_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n440_), .A2(new_n431_), .A3(new_n441_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n443_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n387_), .B2(new_n345_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G226gat), .A2(G233gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT19), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n334_), .B1(KEYINPUT24), .B2(new_n335_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT25), .B(G183gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT87), .ZN(new_n459_));
  INV_X1    g258(.A(new_n329_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n336_), .A2(KEYINPUT24), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT88), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n335_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n342_), .B(KEYINPUT89), .ZN(new_n465_));
  INV_X1    g264(.A(G176gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n334_), .B1(G183gat), .B2(G190gat), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n468_), .A2(new_n336_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n461_), .A2(new_n464_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n416_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n453_), .A2(new_n456_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT90), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n387_), .A2(new_n470_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n345_), .A2(new_n416_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n452_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n473_), .B1(new_n476_), .B2(new_n456_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n476_), .A2(new_n473_), .A3(new_n456_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n472_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G8gat), .B(G36gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT18), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G64gat), .B(G92gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n472_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n476_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(KEYINPUT90), .A3(new_n455_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n489_), .B2(new_n477_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n484_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT27), .B1(new_n486_), .B2(new_n491_), .ZN(new_n492_));
  AOI211_X1 g291(.A(new_n487_), .B(new_n485_), .C1(new_n489_), .C2(new_n477_), .ZN(new_n493_));
  AOI211_X1 g292(.A(new_n452_), .B(new_n455_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n418_), .A2(new_n419_), .A3(new_n470_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n456_), .B1(new_n495_), .B2(new_n453_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT27), .B1(new_n497_), .B2(new_n484_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n413_), .A2(KEYINPUT91), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n407_), .A2(new_n501_), .A3(new_n412_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n502_), .A3(new_n363_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(new_n363_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT92), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n445_), .A2(new_n510_), .A3(new_n413_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n507_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n509_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G29gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT0), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(new_n300_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G85gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n509_), .B(new_n518_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n492_), .A2(new_n499_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n512_), .A2(new_n508_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n511_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n518_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n521_), .A2(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n486_), .A2(new_n491_), .A3(new_n525_), .A4(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n494_), .A2(new_n496_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n484_), .A2(KEYINPUT32), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT94), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n532_), .B(KEYINPUT93), .Z(new_n535_));
  NAND2_X1  g334(.A1(new_n490_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n537_), .A3(new_n532_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n534_), .A2(new_n536_), .A3(new_n522_), .A4(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n530_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n372_), .B1(new_n449_), .B2(new_n448_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n451_), .A2(new_n523_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n305_), .B(new_n230_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT65), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n240_), .A2(new_n306_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT64), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n306_), .A2(KEYINPUT12), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n255_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n543_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n545_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n550_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n550_), .A2(new_n558_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(KEYINPUT13), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT13), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n243_), .A2(new_n291_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n212_), .A2(new_n291_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n212_), .B(new_n291_), .Z(new_n576_));
  INV_X1    g375(.A(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G169gat), .B(G197gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT75), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT74), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n581_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n579_), .B(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n570_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n542_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n321_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT95), .Z(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n286_), .A3(new_n522_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT38), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n587_), .A2(new_n319_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT96), .Z(new_n595_));
  NOR2_X1   g394(.A1(new_n272_), .A2(new_n276_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n542_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n522_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G1gat), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n593_), .A2(new_n600_), .ZN(G1324gat));
  NOR2_X1   g400(.A1(new_n492_), .A2(new_n499_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n591_), .A2(new_n287_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G8gat), .B1(new_n598_), .B2(new_n602_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT39), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(G1325gat));
  OAI21_X1  g408(.A(G15gat), .B1(new_n598_), .B2(new_n447_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT41), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n591_), .A2(new_n352_), .A3(new_n372_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1326gat));
  INV_X1    g412(.A(G22gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n448_), .A2(new_n449_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n591_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G22gat), .B1(new_n598_), .B2(new_n615_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT97), .B(KEYINPUT42), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(G1327gat));
  OAI21_X1  g420(.A(KEYINPUT43), .B1(new_n542_), .B2(new_n284_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n277_), .A2(new_n283_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT27), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n490_), .A2(new_n484_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n626_), .B2(new_n493_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n493_), .A2(new_n498_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n599_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n450_), .B2(new_n443_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n541_), .A2(new_n540_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n623_), .B(new_n624_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n319_), .B1(new_n622_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(new_n587_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT44), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(G29gat), .A3(new_n522_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(KEYINPUT44), .ZN(new_n637_));
  INV_X1    g436(.A(new_n596_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n319_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n589_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n599_), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n636_), .A2(new_n637_), .B1(G29gat), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1328gat));
  INV_X1    g443(.A(G36gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n637_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n602_), .B1(new_n634_), .B2(KEYINPUT44), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n640_), .A2(G36gat), .A3(new_n602_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT99), .B(KEYINPUT45), .Z(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n654_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n649_), .A2(new_n656_), .A3(new_n658_), .A4(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n656_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n662_), .B2(new_n648_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1329gat));
  OAI21_X1  g463(.A(new_n349_), .B1(new_n640_), .B2(new_n447_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n635_), .A2(G43gat), .A3(new_n372_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n637_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g467(.A1(new_n640_), .A2(new_n615_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(G50gat), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n635_), .A2(G50gat), .A3(new_n616_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n646_), .ZN(G1331gat));
  XNOR2_X1  g471(.A(new_n579_), .B(new_n584_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n570_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n542_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n321_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n300_), .A3(new_n522_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n674_), .A2(new_n673_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n597_), .A2(new_n319_), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n599_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(G1332gat));
  OAI21_X1  g480(.A(G64gat), .B1(new_n679_), .B2(new_n602_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT103), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT102), .B(KEYINPUT48), .Z(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n684_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n603_), .A2(new_n298_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT104), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n676_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n686_), .A3(new_n689_), .ZN(G1333gat));
  OAI21_X1  g489(.A(G71gat), .B1(new_n679_), .B2(new_n447_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT49), .ZN(new_n692_));
  INV_X1    g491(.A(G71gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n676_), .A2(new_n693_), .A3(new_n372_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1334gat));
  OAI21_X1  g494(.A(G78gat), .B1(new_n679_), .B2(new_n615_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(G78gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n676_), .A2(new_n699_), .A3(new_n616_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1335gat));
  AND2_X1   g500(.A1(new_n675_), .A2(new_n639_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n225_), .A3(new_n522_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n622_), .A2(new_n632_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n319_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n678_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n633_), .A2(KEYINPUT106), .A3(new_n678_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n599_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n703_), .B1(new_n710_), .B2(new_n225_), .ZN(G1336gat));
  NAND3_X1  g510(.A1(new_n702_), .A2(new_n226_), .A3(new_n603_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n602_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n226_), .ZN(G1337gat));
  NAND4_X1  g513(.A1(new_n702_), .A2(new_n221_), .A3(new_n223_), .A4(new_n372_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n447_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n232_), .ZN(new_n718_));
  AND4_X1   g517(.A1(KEYINPUT106), .A2(new_n704_), .A3(new_n705_), .A4(new_n678_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT106), .B1(new_n633_), .B2(new_n678_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n372_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n721_), .B2(G99gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n715_), .B1(new_n718_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT51), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n715_), .C1(new_n718_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1338gat));
  NAND3_X1  g526(.A1(new_n702_), .A2(new_n222_), .A3(new_n616_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n633_), .A2(new_n616_), .A3(new_n678_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G106gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G106gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g533(.A(new_n673_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n277_), .A2(new_n283_), .A3(new_n319_), .A4(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n736_), .B(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n673_), .A2(new_n566_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT65), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n543_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n554_), .A2(KEYINPUT65), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n553_), .A2(new_n743_), .A3(new_n744_), .A4(new_n557_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n549_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(KEYINPUT109), .A3(new_n549_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n558_), .A2(KEYINPUT55), .ZN(new_n751_));
  AOI22_X1  g550(.A1(new_n255_), .A2(new_n552_), .B1(new_n545_), .B2(new_n556_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n555_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n741_), .B1(new_n750_), .B2(new_n755_), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n747_), .B(new_n548_), .C1(new_n752_), .C2(new_n544_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT109), .B1(new_n745_), .B2(new_n549_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n741_), .B(new_n755_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n563_), .B1(new_n756_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT110), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n759_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(KEYINPUT56), .A3(new_n563_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n740_), .B1(new_n763_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n579_), .A2(new_n584_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n585_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(KEYINPUT111), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(KEYINPUT111), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n574_), .B2(new_n573_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n567_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n638_), .B1(new_n768_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n566_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n586_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT56), .B1(new_n766_), .B2(new_n563_), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n762_), .B(new_n565_), .C1(new_n765_), .C2(new_n759_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n776_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(KEYINPUT57), .A3(new_n638_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n774_), .A2(new_n780_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT58), .B(new_n788_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n624_), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n779_), .A2(new_n787_), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n739_), .B1(new_n794_), .B2(new_n705_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n603_), .A2(new_n599_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n372_), .A3(new_n615_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT59), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n624_), .A2(new_n792_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n763_), .A2(new_n767_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT58), .B1(new_n800_), .B2(new_n788_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT57), .B1(new_n786_), .B2(new_n638_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT112), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n779_), .A2(new_n805_), .A3(new_n793_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n787_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n739_), .B1(new_n807_), .B2(new_n705_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n797_), .A2(KEYINPUT59), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n798_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT113), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n798_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n586_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n795_), .A2(new_n797_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n815_), .B1(new_n819_), .B2(new_n586_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n817_), .A2(KEYINPUT114), .A3(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1340gat));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n674_), .B2(KEYINPUT60), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT115), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n818_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n826_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT116), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n811_), .A2(new_n674_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n832_), .B2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n818_), .B2(new_n319_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT117), .Z(new_n835_));
  AND2_X1   g634(.A1(new_n812_), .A2(new_n814_), .ZN(new_n836_));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n705_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n835_), .B1(new_n836_), .B2(new_n838_), .ZN(G1342gat));
  NAND3_X1  g638(.A1(new_n812_), .A2(new_n624_), .A3(new_n814_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G134gat), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n638_), .A2(G134gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n819_), .B2(new_n842_), .ZN(G1343gat));
  INV_X1    g642(.A(new_n795_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n603_), .A2(new_n450_), .A3(new_n599_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT118), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n586_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(new_n396_), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n674_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT119), .B(G148gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1345gat));
  NOR2_X1   g651(.A1(new_n847_), .A2(new_n705_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT61), .B(G155gat), .Z(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1346gat));
  OAI21_X1  g654(.A(G162gat), .B1(new_n847_), .B2(new_n284_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n638_), .A2(G162gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n847_), .B2(new_n857_), .ZN(G1347gat));
  NOR2_X1   g657(.A1(new_n447_), .A2(new_n522_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n603_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n616_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n787_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n779_), .A2(new_n793_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(KEYINPUT112), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n319_), .B1(new_n864_), .B2(new_n806_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n673_), .B(new_n861_), .C1(new_n865_), .C2(new_n739_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G169gat), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n861_), .B1(new_n865_), .B2(new_n739_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n673_), .A3(new_n465_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n870_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT120), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n869_), .A2(new_n873_), .A3(new_n876_), .A4(new_n870_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n872_), .B2(new_n570_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n795_), .A2(new_n616_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n603_), .A2(new_n570_), .A3(G176gat), .A4(new_n859_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n879_), .B1(new_n880_), .B2(new_n882_), .ZN(G1349gat));
  NOR3_X1   g682(.A1(new_n871_), .A2(new_n705_), .A3(new_n459_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n880_), .A2(new_n319_), .A3(new_n603_), .A4(new_n859_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n330_), .B2(new_n885_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n871_), .B2(new_n284_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n596_), .A2(new_n460_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT121), .Z(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n871_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1351gat));
  NOR3_X1   g691(.A1(new_n602_), .A2(new_n522_), .A3(new_n450_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n795_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n673_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n381_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT124), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n899_), .A3(new_n381_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n895_), .A2(G197gat), .A3(new_n673_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n903_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT125), .B1(new_n901_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n898_), .A2(new_n900_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n908_), .A2(new_n909_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(G1352gat));
  NAND2_X1  g710(.A1(new_n895_), .A2(new_n570_), .ZN(new_n912_));
  XOR2_X1   g711(.A(KEYINPUT126), .B(G204gat), .Z(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1353gat));
  INV_X1    g713(.A(new_n895_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n319_), .A2(new_n916_), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT127), .Z(new_n918_));
  NOR2_X1   g717(.A1(new_n915_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1354gat));
  OR3_X1    g720(.A1(new_n915_), .A2(G218gat), .A3(new_n638_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G218gat), .B1(new_n915_), .B2(new_n284_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1355gat));
endmodule


