//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_;
  XOR2_X1   g000(.A(KEYINPUT22), .B(G169gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT83), .B(G176gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT23), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(G183gat), .B2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT82), .Z(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT26), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n214_), .A2(G190gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n214_), .A2(G190gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n217_), .A2(KEYINPUT79), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(KEYINPUT79), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT80), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT81), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n206_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n224_), .A2(new_n225_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(new_n209_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n211_), .B1(new_n222_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G197gat), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n231_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(G204gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT91), .B1(new_n231_), .B2(G204gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT93), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n236_), .A2(KEYINPUT21), .A3(new_n239_), .A4(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n231_), .A2(G204gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT21), .B1(new_n242_), .B2(new_n233_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n237_), .B(new_n243_), .C1(new_n235_), .C2(KEYINPUT21), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT20), .B1(new_n230_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G226gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT19), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n228_), .A2(new_n208_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n223_), .A2(new_n225_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n206_), .A2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n215_), .A2(new_n217_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT95), .Z(new_n253_));
  OAI211_X1 g052(.A(new_n249_), .B(new_n251_), .C1(new_n253_), .C2(new_n213_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n210_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n241_), .A2(new_n244_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n246_), .A2(new_n248_), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259_));
  INV_X1    g058(.A(G92gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT18), .B(G64gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n230_), .A2(new_n245_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(new_n256_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(KEYINPUT20), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n248_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n258_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n248_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n266_), .A2(KEYINPUT20), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n265_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n246_), .A2(new_n248_), .A3(new_n257_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n263_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n248_), .B1(new_n246_), .B2(new_n257_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n248_), .B2(new_n267_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n263_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(KEYINPUT27), .A3(new_n269_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G22gat), .B(G50gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(G155gat), .B2(G162gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n289_), .A2(KEYINPUT3), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT2), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(KEYINPUT3), .B2(new_n289_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n286_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n287_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT1), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n295_), .B(new_n291_), .C1(new_n285_), .C2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT29), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n300_), .A2(new_n301_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n282_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n304_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n282_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n302_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(KEYINPUT29), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n256_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G228gat), .ZN(new_n312_));
  INV_X1    g111(.A(G233gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT94), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n256_), .B(new_n310_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n309_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G78gat), .B(G106gat), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n321_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n323_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n277_), .B(new_n281_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G57gat), .B(G85gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335_));
  INV_X1    g134(.A(G120gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT86), .B(G113gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n299_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n299_), .A2(new_n339_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(KEYINPUT4), .A3(new_n341_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n341_), .A2(KEYINPUT4), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n343_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n334_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n345_), .A2(new_n348_), .A3(new_n334_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT100), .B1(new_n328_), .B2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n277_), .A2(new_n281_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n327_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n325_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT100), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .A4(new_n352_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n326_), .A2(new_n327_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n258_), .A2(new_n268_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n362_));
  OAI22_X1  g161(.A1(new_n350_), .A2(new_n351_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT98), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n279_), .A2(new_n364_), .A3(new_n362_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n279_), .B2(new_n362_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n363_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT33), .B(new_n334_), .C1(new_n345_), .C2(new_n348_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT97), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT33), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n349_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n342_), .A2(new_n344_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n346_), .A2(new_n343_), .A3(new_n347_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n333_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n371_), .A2(new_n269_), .A3(new_n274_), .A4(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n369_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n360_), .B1(new_n367_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n354_), .A2(new_n359_), .A3(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G15gat), .B(G43gat), .Z(new_n379_));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n384_), .A2(KEYINPUT84), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(KEYINPUT84), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT85), .B1(new_n339_), .B2(KEYINPUT31), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(KEYINPUT31), .B2(new_n339_), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(KEYINPUT87), .Z(new_n390_));
  AND2_X1   g189(.A1(new_n386_), .A2(new_n383_), .ZN(new_n391_));
  OR3_X1    g190(.A1(new_n387_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n387_), .B2(new_n391_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n378_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT101), .ZN(new_n397_));
  INV_X1    g196(.A(new_n355_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(new_n357_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n394_), .A3(new_n352_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT101), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n378_), .A2(new_n401_), .A3(new_n395_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT13), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT70), .B(KEYINPUT5), .Z(new_n405_));
  XNOR2_X1  g204(.A(G120gat), .B(G148gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G176gat), .B(G204gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT10), .B(G99gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(G106gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT64), .ZN(new_n413_));
  AND3_X1   g212(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G85gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n260_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G85gat), .A2(G92gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT9), .A3(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n416_), .B(new_n420_), .C1(KEYINPUT9), .C2(new_n419_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n413_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT7), .ZN(new_n424_));
  INV_X1    g223(.A(G99gat), .ZN(new_n425_));
  INV_X1    g224(.A(G106gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G99gat), .A2(G106gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n427_), .A2(new_n430_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT65), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT66), .ZN(new_n435_));
  AND2_X1   g234(.A1(G85gat), .A2(G92gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n418_), .A2(KEYINPUT66), .A3(new_n419_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT8), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT65), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n416_), .A2(new_n441_), .A3(new_n432_), .A4(new_n427_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n434_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT67), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n434_), .A2(new_n440_), .A3(new_n442_), .A4(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT8), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n438_), .A2(new_n439_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n433_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT68), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n453_));
  AOI211_X1 g252(.A(new_n453_), .B(new_n450_), .C1(new_n444_), .C2(new_n446_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n423_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G57gat), .B(G64gat), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n458_));
  XOR2_X1   g257(.A(G71gat), .B(G78gat), .Z(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n455_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n450_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n462_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n466_), .A2(new_n422_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n466_), .B2(new_n422_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G230gat), .A2(G233gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n465_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT69), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT69), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n465_), .A2(new_n470_), .A3(new_n474_), .A4(new_n471_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n468_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n471_), .B1(new_n477_), .B2(new_n469_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n410_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n409_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n404_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n480_), .A2(new_n409_), .ZN(new_n483_));
  AOI211_X1 g282(.A(new_n478_), .B(new_n410_), .C1(new_n473_), .C2(new_n475_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n483_), .A2(new_n484_), .A3(KEYINPUT13), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT75), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(G1gat), .B2(G8gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT76), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G1gat), .B(G8gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G29gat), .B(G36gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G43gat), .B(G50gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT15), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n497_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n494_), .A2(new_n497_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT78), .A3(new_n502_), .ZN(new_n505_));
  OR3_X1    g304(.A1(new_n494_), .A2(KEYINPUT78), .A3(new_n497_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n503_), .B1(new_n507_), .B2(new_n501_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G169gat), .B(G197gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n508_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n486_), .A2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n403_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n455_), .A2(new_n498_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT34), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n466_), .A2(new_n422_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n524_), .A2(new_n497_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n516_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n516_), .B2(new_n525_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G134gat), .B(G162gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT36), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT72), .B1(new_n528_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n447_), .A2(new_n451_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n453_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n466_), .A2(KEYINPUT68), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n422_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n525_), .B1(new_n538_), .B2(new_n499_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n522_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n516_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n540_), .A2(KEYINPUT72), .A3(new_n533_), .A4(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT73), .B1(new_n534_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n533_), .A3(new_n541_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT72), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n542_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n531_), .B(KEYINPUT36), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT37), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n544_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n547_), .A2(new_n542_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(KEYINPUT74), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n540_), .A2(new_n541_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT74), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(new_n550_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n555_), .B1(new_n556_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n494_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n467_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G211gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT16), .B(G183gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT17), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n569_), .A2(KEYINPUT17), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n554_), .A2(new_n562_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT77), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n515_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n352_), .A2(G1gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT103), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT103), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n579_), .A2(new_n584_), .A3(KEYINPUT38), .A4(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n547_), .A2(new_n542_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n574_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n515_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G1gat), .B1(new_n591_), .B2(new_n352_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT38), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n581_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n585_), .A3(new_n594_), .ZN(G1324gat));
  XNOR2_X1  g394(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G8gat), .B1(new_n591_), .B2(new_n355_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n515_), .A2(KEYINPUT102), .A3(new_n576_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n577_), .A2(new_n578_), .ZN(new_n602_));
  AOI211_X1 g401(.A(G8gat), .B(new_n355_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n597_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n598_), .B(KEYINPUT39), .ZN(new_n605_));
  INV_X1    g404(.A(G8gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n579_), .A2(new_n606_), .A3(new_n398_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n607_), .A3(new_n596_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n604_), .A2(new_n608_), .ZN(G1325gat));
  OAI21_X1  g408(.A(G15gat), .B1(new_n591_), .B2(new_n395_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT41), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT41), .ZN(new_n612_));
  OR3_X1    g411(.A1(new_n577_), .A2(G15gat), .A3(new_n395_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(G1326gat));
  OAI21_X1  g413(.A(G22gat), .B1(new_n591_), .B2(new_n360_), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  OR3_X1    g417(.A1(new_n577_), .A2(G22gat), .A3(new_n360_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(G1327gat));
  NAND2_X1  g419(.A1(new_n554_), .A2(new_n562_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n402_), .A2(new_n400_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n401_), .B1(new_n378_), .B2(new_n395_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n625_));
  NAND2_X1  g424(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n403_), .A2(KEYINPUT106), .A3(KEYINPUT43), .A4(new_n621_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n486_), .A2(new_n513_), .A3(new_n574_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n627_), .A2(new_n628_), .A3(KEYINPUT44), .A4(new_n629_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n353_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G29gat), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n587_), .A2(new_n574_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n403_), .A2(new_n514_), .A3(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n352_), .A2(G29gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n635_), .B1(new_n637_), .B2(new_n638_), .ZN(G1328gat));
  NAND3_X1  g438(.A1(new_n632_), .A2(new_n398_), .A3(new_n633_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G36gat), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n355_), .A2(G36gat), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n515_), .A2(new_n642_), .A3(new_n636_), .A4(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n643_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT107), .B1(new_n637_), .B2(new_n645_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n644_), .A2(KEYINPUT45), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT45), .B1(new_n644_), .B2(new_n646_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n641_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n641_), .A2(new_n649_), .A3(KEYINPUT46), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NAND3_X1  g453(.A1(new_n632_), .A2(new_n394_), .A3(new_n633_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G43gat), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n637_), .A2(G43gat), .A3(new_n395_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT47), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(KEYINPUT47), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1330gat));
  OR3_X1    g461(.A1(new_n637_), .A2(G50gat), .A3(new_n360_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n632_), .A2(new_n357_), .A3(new_n633_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G50gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G50gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(G1331gat));
  AND3_X1   g467(.A1(new_n403_), .A2(new_n513_), .A3(new_n486_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(new_n576_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G57gat), .B1(new_n670_), .B2(new_n353_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n590_), .ZN(new_n672_));
  INV_X1    g471(.A(G57gat), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n352_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n671_), .A2(new_n674_), .ZN(G1332gat));
  OAI21_X1  g474(.A(G64gat), .B1(new_n672_), .B2(new_n355_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT48), .ZN(new_n677_));
  INV_X1    g476(.A(G64gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n670_), .A2(new_n678_), .A3(new_n398_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1333gat));
  OAI21_X1  g479(.A(G71gat), .B1(new_n672_), .B2(new_n395_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT49), .ZN(new_n682_));
  INV_X1    g481(.A(G71gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n670_), .A2(new_n683_), .A3(new_n394_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1334gat));
  OAI21_X1  g484(.A(G78gat), .B1(new_n672_), .B2(new_n360_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT50), .ZN(new_n687_));
  INV_X1    g486(.A(G78gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n670_), .A2(new_n688_), .A3(new_n357_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1335gat));
  NAND2_X1  g489(.A1(new_n669_), .A2(new_n636_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n417_), .B1(new_n691_), .B2(new_n352_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n486_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(new_n512_), .A3(new_n574_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n352_), .A2(new_n417_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT109), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n627_), .A2(new_n628_), .A3(new_n694_), .A4(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n692_), .A2(new_n697_), .ZN(G1336gat));
  OAI21_X1  g497(.A(new_n260_), .B1(new_n691_), .B2(new_n355_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n355_), .A2(new_n260_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n627_), .A2(new_n628_), .A3(new_n694_), .A4(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n699_), .A2(new_n700_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n701_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n701_), .A2(KEYINPUT111), .A3(new_n703_), .A4(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1337gat));
  AND4_X1   g508(.A1(new_n394_), .A2(new_n627_), .A3(new_n628_), .A4(new_n694_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n395_), .A2(new_n411_), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n710_), .A2(new_n425_), .B1(new_n691_), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g512(.A1(new_n627_), .A2(new_n628_), .A3(new_n357_), .A4(new_n694_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(G106gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G106gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n357_), .A2(new_n426_), .ZN(new_n718_));
  OAI22_X1  g517(.A1(new_n716_), .A2(new_n717_), .B1(new_n691_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT53), .ZN(G1339gat));
  OR2_X1    g519(.A1(new_n508_), .A2(new_n511_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n505_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n500_), .A2(new_n502_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n722_), .B(new_n511_), .C1(new_n501_), .C2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(new_n484_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n473_), .A2(new_n475_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT55), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n465_), .A2(new_n470_), .A3(KEYINPUT55), .A4(new_n471_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n465_), .A2(new_n470_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n471_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT56), .B1(new_n734_), .B2(new_n410_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT55), .B1(new_n473_), .B2(new_n475_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT56), .B(new_n410_), .C1(new_n736_), .C2(new_n732_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT58), .B(new_n726_), .C1(new_n735_), .C2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n410_), .B1(new_n736_), .B2(new_n732_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT56), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n737_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n726_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT58), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n745_), .A2(KEYINPUT114), .A3(KEYINPUT58), .A4(new_n726_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n741_), .A2(new_n748_), .A3(new_n621_), .A4(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n725_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n744_), .A2(KEYINPUT113), .A3(new_n737_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n512_), .B(new_n481_), .C1(new_n737_), .C2(KEYINPUT113), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(KEYINPUT57), .A3(new_n587_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n481_), .A2(new_n512_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n738_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n744_), .A2(KEYINPUT113), .A3(new_n737_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n751_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n762_), .B2(new_n588_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n750_), .A2(new_n756_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n589_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n513_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT112), .B1(new_n575_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n552_), .B1(new_n586_), .B2(KEYINPUT73), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n549_), .A2(new_n768_), .B1(new_n587_), .B2(new_n555_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n479_), .A2(new_n404_), .A3(new_n481_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT13), .B1(new_n483_), .B2(new_n484_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n512_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n769_), .A2(new_n770_), .A3(new_n773_), .A4(new_n574_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n767_), .A2(KEYINPUT54), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT54), .B1(new_n767_), .B2(new_n774_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n352_), .B1(new_n765_), .B2(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n395_), .A2(new_n357_), .A3(new_n398_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT59), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n782_), .B2(KEYINPUT59), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n783_), .ZN(new_n786_));
  INV_X1    g585(.A(G113gat), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n513_), .A2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n780_), .A2(KEYINPUT115), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n780_), .A2(KEYINPUT115), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n512_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n786_), .A2(new_n788_), .B1(new_n791_), .B2(new_n787_), .ZN(G1340gat));
  NAND2_X1  g591(.A1(new_n785_), .A2(new_n783_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(new_n486_), .C1(new_n781_), .C2(new_n783_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G120gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n336_), .B1(new_n693_), .B2(KEYINPUT60), .ZN(new_n796_));
  OAI221_X1 g595(.A(new_n796_), .B1(KEYINPUT60), .B2(new_n336_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1341gat));
  INV_X1    g597(.A(G127gat), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n589_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n574_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n786_), .A2(new_n800_), .B1(new_n801_), .B2(new_n799_), .ZN(G1342gat));
  NAND2_X1  g601(.A1(new_n621_), .A2(G134gat), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT117), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n588_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n805_));
  INV_X1    g604(.A(G134gat), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n786_), .A2(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(G1343gat));
  NOR2_X1   g606(.A1(new_n394_), .A2(new_n328_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n764_), .A2(new_n589_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n776_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n767_), .A2(new_n774_), .A3(KEYINPUT54), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n353_), .B(new_n808_), .C1(new_n809_), .C2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT118), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n778_), .A2(new_n815_), .A3(new_n808_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n512_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n486_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n574_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT119), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n817_), .A2(new_n824_), .A3(new_n574_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT61), .B(G155gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n826_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n824_), .B1(new_n817_), .B2(new_n574_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT119), .B(new_n589_), .C1(new_n814_), .C2(new_n816_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(G1346gat));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n765_), .A2(new_n777_), .ZN(new_n834_));
  AND4_X1   g633(.A1(new_n815_), .A2(new_n834_), .A3(new_n353_), .A4(new_n808_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n815_), .B1(new_n778_), .B2(new_n808_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n621_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G162gat), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n587_), .A2(G162gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n833_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n769_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n842_));
  INV_X1    g641(.A(G162gat), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n833_), .B(new_n840_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n841_), .A2(new_n845_), .ZN(G1347gat));
  INV_X1    g645(.A(G169gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n357_), .B1(new_n765_), .B2(new_n777_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n395_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n512_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(KEYINPUT121), .Z(new_n851_));
  AOI21_X1  g650(.A(new_n847_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT62), .Z(new_n853_));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n849_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT122), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n513_), .A2(new_n202_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n853_), .B1(new_n855_), .B2(new_n856_), .ZN(G1348gat));
  INV_X1    g656(.A(new_n855_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n203_), .B1(new_n858_), .B2(new_n486_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n854_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n860_), .A2(G176gat), .A3(new_n486_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1349gat));
  AOI21_X1  g661(.A(G183gat), .B1(new_n860_), .B2(new_n574_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n589_), .A2(new_n212_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n858_), .B2(new_n864_), .ZN(G1350gat));
  OAI21_X1  g664(.A(G190gat), .B1(new_n855_), .B2(new_n769_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n587_), .A2(new_n253_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n855_), .B2(new_n867_), .ZN(G1351gat));
  NAND4_X1  g667(.A1(new_n395_), .A2(new_n352_), .A3(new_n398_), .A4(new_n357_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n765_), .B2(new_n777_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n512_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n231_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(KEYINPUT123), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n872_), .A2(KEYINPUT123), .ZN(new_n874_));
  AOI211_X1 g673(.A(new_n873_), .B(new_n874_), .C1(new_n231_), .C2(new_n871_), .ZN(G1352gat));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n486_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n870_), .A2(KEYINPUT124), .A3(new_n486_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(G204gat), .A3(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n876_), .A2(G204gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(KEYINPUT125), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(KEYINPUT125), .B2(new_n880_), .ZN(G1353gat));
  NAND2_X1  g682(.A1(new_n870_), .A2(new_n574_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  AND2_X1   g684(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n884_), .B2(new_n885_), .ZN(G1354gat));
  INV_X1    g687(.A(G218gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n870_), .A2(new_n889_), .A3(new_n588_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n870_), .A2(new_n621_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(KEYINPUT126), .Z(G1355gat));
endmodule


