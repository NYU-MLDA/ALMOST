//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  AND3_X1   g002(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(KEYINPUT78), .B1(G183gat), .B2(G190gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT77), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT77), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n210_));
  AND2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI22_X1  g011(.A1(KEYINPUT23), .A2(new_n206_), .B1(new_n212_), .B2(KEYINPUT81), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT81), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(new_n211_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n203_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT79), .B(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT22), .B(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT80), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n218_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n206_), .A2(KEYINPUT23), .B1(new_n214_), .B2(new_n211_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT75), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  INV_X1    g026(.A(G176gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT24), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G183gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT74), .B1(new_n233_), .B2(KEYINPUT25), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n234_), .B(new_n235_), .C1(new_n236_), .C2(KEYINPUT74), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n225_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n229_), .A2(new_n230_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(KEYINPUT76), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n229_), .A2(new_n230_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(new_n240_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  OAI22_X1  g045(.A1(new_n217_), .A2(new_n224_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT30), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT83), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G15gat), .B(G43gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G71gat), .B(G99gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n253_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n218_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n223_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n206_), .A2(KEYINPUT23), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n212_), .A2(KEYINPUT81), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n216_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n203_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n237_), .A2(new_n232_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n268_), .A2(new_n225_), .A3(new_n245_), .A4(new_n242_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n269_), .A3(KEYINPUT30), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n249_), .A2(new_n257_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT84), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n249_), .A2(new_n270_), .A3(KEYINPUT84), .A4(new_n257_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n257_), .B1(new_n249_), .B2(new_n270_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT31), .ZN(new_n279_));
  XOR2_X1   g078(.A(G127gat), .B(G134gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(G113gat), .B(G120gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G113gat), .B(G120gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT85), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n282_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n275_), .A2(new_n290_), .A3(new_n277_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n279_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n289_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n290_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n294_));
  AOI211_X1 g093(.A(KEYINPUT31), .B(new_n276_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(G141gat), .ZN(new_n300_));
  INV_X1    g099(.A(G148gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT1), .ZN(new_n304_));
  OR2_X1    g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n303_), .A2(KEYINPUT1), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n299_), .B(new_n302_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT3), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n299_), .A2(KEYINPUT2), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n299_), .A2(KEYINPUT2), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n310_), .A2(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n303_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n308_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n316_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT28), .B1(new_n316_), .B2(KEYINPUT29), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G22gat), .B(G50gat), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G78gat), .B(G106gat), .ZN(new_n323_));
  AND2_X1   g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT86), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT21), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n330_), .B(new_n331_), .C1(new_n328_), .C2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n328_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n331_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n332_), .A4(KEYINPUT21), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n326_), .B1(new_n327_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n324_), .A2(new_n325_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n327_), .A2(new_n325_), .A3(new_n338_), .A4(new_n324_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n323_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n322_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n342_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n323_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n341_), .A2(new_n342_), .A3(new_n323_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n345_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT20), .ZN(new_n352_));
  INV_X1    g151(.A(new_n338_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n247_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT23), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n211_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n265_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n258_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n264_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n244_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n236_), .A2(new_n235_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n365_), .A2(new_n258_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n366_), .B(new_n367_), .C1(new_n368_), .C2(new_n244_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n338_), .B(new_n363_), .C1(new_n364_), .C2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n352_), .B1(new_n354_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT90), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT19), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n338_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n370_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT20), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT90), .B1(new_n379_), .B2(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n247_), .A2(new_n338_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT20), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n363_), .B1(new_n364_), .B2(new_n369_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n375_), .B1(new_n383_), .B2(new_n338_), .ZN(new_n384_));
  OAI22_X1  g183(.A1(new_n376_), .A2(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  XOR2_X1   g185(.A(G64gat), .B(G92gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G8gat), .B(G36gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT92), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n389_), .B(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(new_n386_), .A3(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n382_), .A2(new_n384_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n372_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n379_), .A2(KEYINPUT90), .A3(new_n374_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n392_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT93), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n397_), .A2(new_n398_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n393_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT94), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT94), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n393_), .B(new_n403_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n316_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n310_), .A2(new_n311_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n312_), .A2(new_n313_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n303_), .B(new_n305_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n282_), .A2(new_n285_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n308_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT0), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT97), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G57gat), .B(G85gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n405_), .A2(new_n410_), .A3(KEYINPUT4), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT95), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n405_), .A2(new_n410_), .A3(KEYINPUT95), .A4(KEYINPUT4), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT96), .B(KEYINPUT4), .Z(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n408_), .B2(new_n308_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n289_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(new_n412_), .ZN(new_n429_));
  AOI211_X1 g228(.A(new_n414_), .B(new_n420_), .C1(new_n425_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n420_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n411_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n413_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n428_), .A2(new_n413_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n425_), .A2(new_n434_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n430_), .A2(KEYINPUT33), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n430_), .A2(new_n437_), .A3(KEYINPUT33), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n425_), .A2(new_n429_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n414_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n431_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT98), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n436_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n402_), .A2(new_n404_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n430_), .A2(KEYINPUT100), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT100), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n441_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n414_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n447_), .B(new_n449_), .C1(new_n450_), .C2(new_n431_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n397_), .B1(new_n452_), .B2(new_n392_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n383_), .A2(KEYINPUT99), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n383_), .A2(KEYINPUT99), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n338_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n374_), .B1(new_n456_), .B2(new_n382_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(KEYINPUT32), .A3(new_n398_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(new_n453_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n351_), .B1(new_n446_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT27), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n397_), .A2(new_n398_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n458_), .B2(new_n392_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n401_), .A2(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n351_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(new_n451_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n298_), .B1(new_n461_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n401_), .A2(new_n462_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n451_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n351_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n463_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT101), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT101), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n465_), .A2(new_n477_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G120gat), .B(G148gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT5), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G176gat), .B(G204gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT10), .B(G99gat), .Z(new_n486_));
  INV_X1    g285(.A(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G85gat), .B(G92gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n490_));
  INV_X1    g289(.A(G85gat), .ZN(new_n491_));
  INV_X1    g290(.A(G92gat), .ZN(new_n492_));
  OR3_X1    g291(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT9), .ZN(new_n493_));
  NAND3_X1  g292(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n488_), .A2(new_n490_), .A3(new_n493_), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT7), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n496_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT64), .A3(new_n494_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n499_), .B1(new_n506_), .B2(new_n489_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n489_), .A2(new_n499_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n498_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(G71gat), .B(G78gat), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n511_), .A2(new_n513_), .A3(KEYINPUT11), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n513_), .B1(KEYINPUT11), .B2(new_n511_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n510_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT65), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n510_), .A2(new_n517_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n518_), .A2(KEYINPUT65), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G230gat), .A2(G233gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT12), .B1(new_n510_), .B2(new_n517_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n518_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n510_), .A2(KEYINPUT66), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n529_), .B(new_n498_), .C1(new_n507_), .C2(new_n509_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n528_), .A2(KEYINPUT12), .A3(new_n517_), .A4(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n531_), .A3(new_n524_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n485_), .B1(new_n525_), .B2(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n532_), .B(new_n485_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n533_), .A2(KEYINPUT13), .A3(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT13), .B1(new_n533_), .B2(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G29gat), .B(G36gat), .Z(new_n542_));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G29gat), .B(G36gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT67), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G43gat), .B(G50gat), .Z(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n548_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT73), .B(G15gat), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n556_), .A2(G22gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(G22gat), .ZN(new_n558_));
  INV_X1    g357(.A(G8gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G1gat), .B(G8gat), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n562_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n554_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n555_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n553_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n541_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n552_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n571_), .A2(new_n541_), .A3(new_n569_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n573_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n539_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n480_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT34), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n552_), .A2(KEYINPUT15), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n566_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n588_), .A2(new_n528_), .A3(KEYINPUT68), .A4(new_n530_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n585_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n510_), .B2(new_n552_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT69), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(KEYINPUT69), .B(new_n590_), .C1(new_n510_), .C2(new_n552_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n528_), .A2(new_n555_), .A3(new_n567_), .A4(new_n530_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT68), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n586_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n591_), .A2(new_n586_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n596_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n601_), .B2(new_n596_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n600_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT36), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n606_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT72), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n600_), .A2(new_n605_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT71), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT72), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n616_), .A2(new_n607_), .A3(new_n617_), .A4(new_n611_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n610_), .A2(KEYINPUT36), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n600_), .A2(new_n605_), .A3(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n614_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n565_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n517_), .ZN(new_n625_));
  XOR2_X1   g424(.A(G127gat), .B(G155gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT16), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT17), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n629_), .A2(new_n630_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n625_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n625_), .A2(new_n631_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n622_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n581_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n202_), .B1(new_n638_), .B2(new_n451_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT102), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n615_), .A2(new_n611_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(KEYINPUT37), .A3(new_n620_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT37), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n621_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n636_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n581_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n202_), .A3(new_n451_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT38), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n640_), .A2(new_n650_), .ZN(G1324gat));
  INV_X1    g450(.A(new_n465_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n559_), .B1(new_n638_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT39), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n648_), .A2(new_n559_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(KEYINPUT40), .A3(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1325gat));
  NAND2_X1  g459(.A1(new_n638_), .A2(new_n297_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G15gat), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT41), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT41), .ZN(new_n664_));
  INV_X1    g463(.A(G15gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n648_), .A2(new_n665_), .A3(new_n297_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n664_), .A3(new_n666_), .ZN(G1326gat));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n638_), .B2(new_n351_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT42), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n648_), .A2(new_n668_), .A3(new_n351_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n621_), .A2(new_n635_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n581_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n451_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n645_), .B1(new_n470_), .B2(new_n479_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(KEYINPUT103), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n476_), .A2(new_n478_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n460_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n444_), .B1(new_n401_), .B2(KEYINPUT94), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n404_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n468_), .B1(new_n683_), .B2(new_n351_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n680_), .B1(new_n684_), .B2(new_n298_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n679_), .B(KEYINPUT43), .C1(new_n685_), .C2(new_n645_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n678_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n580_), .A3(new_n636_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(KEYINPUT44), .ZN(new_n690_));
  INV_X1    g489(.A(G29gat), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n472_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(KEYINPUT44), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n675_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n465_), .B1(new_n688_), .B2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n693_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n465_), .B(KEYINPUT104), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n674_), .A2(new_n695_), .A3(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT106), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n698_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n698_), .B2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1329gat));
  AND2_X1   g507(.A1(new_n674_), .A2(new_n297_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(G43gat), .ZN(new_n710_));
  OAI211_X1 g509(.A(G43gat), .B(new_n297_), .C1(new_n689_), .C2(KEYINPUT44), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n688_), .A2(new_n696_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g513(.A(G50gat), .B1(new_n674_), .B2(new_n351_), .ZN(new_n715_));
  INV_X1    g514(.A(G50gat), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n690_), .A2(new_n716_), .A3(new_n466_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n717_), .B2(new_n693_), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n538_), .A2(new_n578_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n480_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n637_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT107), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(G57gat), .A3(new_n451_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT108), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n720_), .A2(new_n647_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n451_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1332gat));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n722_), .B2(new_n700_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT48), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n728_), .A3(new_n700_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n722_), .B2(new_n297_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT49), .Z(new_n735_));
  NAND2_X1  g534(.A1(new_n297_), .A2(new_n733_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT109), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n725_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1334gat));
  INV_X1    g538(.A(G78gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n722_), .B2(new_n351_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT50), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n725_), .A2(new_n740_), .A3(new_n351_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1335gat));
  AND2_X1   g543(.A1(new_n720_), .A2(new_n673_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n491_), .A3(new_n451_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n719_), .A2(new_n636_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n687_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n747_), .B1(new_n678_), .B2(new_n686_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT110), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n472_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n746_), .B1(new_n754_), .B2(new_n491_), .ZN(G1336gat));
  NAND3_X1  g554(.A1(new_n745_), .A2(new_n492_), .A3(new_n652_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n699_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n492_), .ZN(G1337gat));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(KEYINPUT51), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n751_), .A2(new_n753_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n297_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G99gat), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n297_), .A2(new_n486_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n745_), .A2(new_n765_), .B1(new_n759_), .B2(KEYINPUT51), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n761_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n766_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n768_), .B(new_n760_), .C1(new_n763_), .C2(G99gat), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n745_), .A2(new_n487_), .A3(new_n351_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n772_));
  AOI211_X1 g571(.A(new_n466_), .B(new_n747_), .C1(new_n678_), .C2(new_n686_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n487_), .B1(new_n773_), .B2(KEYINPUT112), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT112), .B1(new_n752_), .B2(new_n351_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n772_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n687_), .A2(KEYINPUT112), .A3(new_n351_), .A4(new_n748_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G106gat), .ZN(new_n779_));
  INV_X1    g578(.A(new_n772_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n779_), .A2(new_n775_), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n771_), .B1(new_n777_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n771_), .C1(new_n777_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n532_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n527_), .A2(new_n531_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(G230gat), .A3(G233gat), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n527_), .A2(new_n531_), .A3(KEYINPUT55), .A4(new_n524_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n484_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n484_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n578_), .B(new_n534_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n577_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n568_), .A2(new_n541_), .A3(new_n569_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n571_), .A2(new_n569_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n799_), .B(new_n576_), .C1(new_n800_), .C2(new_n541_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n798_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n621_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n788_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n621_), .A2(new_n804_), .A3(KEYINPUT114), .A4(KEYINPUT57), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n805_), .A2(new_n806_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n802_), .A2(new_n534_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n811_), .B(KEYINPUT58), .C1(new_n795_), .C2(new_n796_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n810_), .B1(new_n645_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n636_), .B1(new_n809_), .B2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n645_), .A2(new_n579_), .A3(new_n538_), .A4(new_n635_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT54), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n465_), .A2(new_n451_), .A3(new_n473_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n823_), .A2(G113gat), .A3(new_n579_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n621_), .A2(new_n644_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n816_), .B1(new_n826_), .B2(new_n642_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT57), .B1(new_n621_), .B2(new_n804_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n810_), .B(new_n830_), .C1(new_n645_), .C2(new_n816_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n807_), .A2(new_n808_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n636_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n833_), .B2(new_n636_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n820_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n822_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n837_), .A2(new_n840_), .B1(new_n823_), .B2(KEYINPUT59), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n841_), .A2(new_n578_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n787_), .B(new_n825_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n841_), .B2(new_n578_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT117), .B1(new_n845_), .B2(new_n824_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(new_n841_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G120gat), .B1(new_n848_), .B2(new_n538_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n823_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n539_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n850_), .A2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT118), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n849_), .A2(new_n856_), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n848_), .B2(new_n636_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n636_), .A2(G127gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n823_), .B2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g659(.A(G134gat), .B1(new_n850_), .B2(new_n622_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n646_), .A2(G134gat), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT119), .Z(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n841_), .B2(new_n863_), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n298_), .A2(new_n351_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n700_), .A2(new_n472_), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n821_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n579_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n300_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n538_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n301_), .ZN(G1345gat));
  NAND3_X1  g670(.A1(new_n821_), .A2(new_n635_), .A3(new_n866_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT120), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  NOR2_X1   g674(.A1(new_n867_), .A2(new_n621_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(G162gat), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n876_), .A2(KEYINPUT121), .A3(G162gat), .ZN(new_n880_));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n867_), .A2(new_n881_), .A3(new_n645_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n879_), .A2(new_n880_), .A3(new_n882_), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n699_), .A2(new_n451_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n297_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n351_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n837_), .A2(new_n578_), .A3(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n837_), .A2(new_n578_), .A3(new_n220_), .A4(new_n886_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT62), .B1(new_n887_), .B2(G169gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT122), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n887_), .A2(G169gat), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n895_), .A2(new_n896_), .A3(new_n888_), .A4(new_n889_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n892_), .A2(new_n897_), .ZN(G1348gat));
  INV_X1    g697(.A(new_n219_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n837_), .A2(new_n886_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n539_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n821_), .A2(new_n466_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT123), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n884_), .A2(G176gat), .A3(new_n539_), .A4(new_n297_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(KEYINPUT124), .A3(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n904_), .A2(new_n905_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n901_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(G1349gat));
  OR3_X1    g710(.A1(new_n904_), .A2(new_n636_), .A3(new_n885_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n636_), .A2(new_n236_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n912_), .A2(new_n233_), .B1(new_n900_), .B2(new_n913_), .ZN(G1350gat));
  INV_X1    g713(.A(new_n900_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G190gat), .B1(new_n915_), .B2(new_n645_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n900_), .A2(new_n235_), .A3(new_n622_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1351gat));
  NOR3_X1   g717(.A1(new_n699_), .A2(new_n451_), .A3(new_n865_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n821_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n578_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g722(.A(G204gat), .ZN(new_n924_));
  OR3_X1    g723(.A1(new_n920_), .A2(KEYINPUT125), .A3(new_n538_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT125), .B1(new_n920_), .B2(new_n538_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT126), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n920_), .A2(new_n538_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n924_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n928_), .B1(new_n927_), .B2(new_n931_), .ZN(G1353gat));
  NAND2_X1  g731(.A1(new_n921_), .A2(new_n635_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  AND2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n936_), .A2(KEYINPUT127), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(KEYINPUT127), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n933_), .A2(new_n934_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .ZN(G1354gat));
  OAI21_X1  g739(.A(G218gat), .B1(new_n920_), .B2(new_n645_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n621_), .A2(G218gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n920_), .B2(new_n942_), .ZN(G1355gat));
endmodule


