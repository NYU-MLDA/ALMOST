//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n968_, new_n969_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1012_, new_n1014_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1025_, new_n1026_;
  INV_X1    g000(.A(KEYINPUT104), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n205_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT9), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT10), .B(G99gat), .Z(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n217_), .A2(new_n218_), .A3(new_n223_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(KEYINPUT66), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT65), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT7), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n230_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n220_), .A2(new_n222_), .A3(new_n236_), .ZN(new_n237_));
  OAI22_X1  g036(.A1(new_n233_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n229_), .A2(new_n235_), .A3(new_n237_), .A4(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n228_), .B1(new_n239_), .B2(new_n211_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n211_), .A2(new_n228_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n235_), .A2(new_n238_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(new_n242_), .B2(new_n223_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n210_), .B(new_n227_), .C1(new_n240_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G230gat), .ZN(new_n245_));
  INV_X1    g044(.A(G233gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n227_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n210_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT12), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n249_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n248_), .B1(new_n252_), .B2(new_n244_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT67), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n250_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n248_), .B(new_n244_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262_));
  INV_X1    g061(.A(new_n257_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G120gat), .B(G148gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G176gat), .B(G204gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n258_), .A2(new_n264_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n261_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT70), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n261_), .A2(new_n263_), .A3(new_n276_), .A4(new_n269_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n258_), .A2(new_n264_), .A3(KEYINPUT69), .A4(new_n270_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n273_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT13), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n273_), .A2(KEYINPUT13), .A3(new_n278_), .A4(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n287_));
  AND4_X1   g086(.A1(new_n217_), .A2(new_n218_), .A3(new_n223_), .A4(new_n226_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n239_), .A2(new_n211_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT8), .ZN(new_n290_));
  INV_X1    g089(.A(new_n243_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n288_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G29gat), .B(G36gat), .Z(new_n293_));
  XOR2_X1   g092(.A(G43gat), .B(G50gat), .Z(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G29gat), .B(G36gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G43gat), .B(G50gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT15), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n298_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT15), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n287_), .B1(new_n292_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G232gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT34), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(KEYINPUT35), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n292_), .B2(new_n301_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n250_), .A2(KEYINPUT73), .A3(new_n300_), .A4(new_n303_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(KEYINPUT35), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT72), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G190gat), .B(G218gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT74), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G134gat), .B(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n317_), .A2(new_n318_), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n320_), .A2(KEYINPUT36), .A3(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n305_), .A2(new_n309_), .A3(new_n310_), .A4(new_n313_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n315_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT36), .B1(new_n320_), .B2(new_n321_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n321_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT36), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n319_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n326_), .A2(new_n329_), .A3(KEYINPUT75), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT75), .B1(new_n326_), .B2(new_n329_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT76), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n329_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(new_n329_), .A3(KEYINPUT75), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n315_), .B2(new_n323_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT37), .B1(new_n325_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT37), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n315_), .A2(new_n323_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n335_), .A2(new_n337_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n342_), .B(new_n324_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n345_), .A3(KEYINPUT77), .ZN(new_n346_));
  OR2_X1    g145(.A1(G1gat), .A2(G8gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G1gat), .A2(G8gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT78), .ZN(new_n350_));
  INV_X1    g149(.A(G15gat), .ZN(new_n351_));
  INV_X1    g150(.A(G22gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G15gat), .A2(G22gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n353_), .A2(new_n354_), .B1(KEYINPUT14), .B2(new_n348_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n347_), .A2(new_n356_), .A3(new_n348_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n350_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n355_), .B1(new_n350_), .B2(new_n357_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G231gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(new_n210_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G127gat), .B(G155gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT16), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G183gat), .B(G211gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT17), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n369_), .A2(KEYINPUT79), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n364_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n369_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n364_), .B(new_n372_), .C1(new_n368_), .C2(new_n370_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n376_), .B(KEYINPUT37), .C1(new_n325_), .C2(new_n340_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n346_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n286_), .A2(KEYINPUT80), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT27), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n383_));
  INV_X1    g182(.A(G204gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(G197gat), .ZN(new_n385_));
  INV_X1    g184(.A(G197gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT21), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(G197gat), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n384_), .A2(G197gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n386_), .A2(G204gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT21), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G211gat), .B(G218gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n385_), .A2(new_n389_), .A3(new_n387_), .ZN(new_n396_));
  INV_X1    g195(.A(G218gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G211gat), .ZN(new_n398_));
  INV_X1    g197(.A(G211gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G218gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n388_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n395_), .A2(KEYINPUT94), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT94), .B1(new_n395_), .B2(new_n402_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G169gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT22), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT22), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G169gat), .ZN(new_n409_));
  INV_X1    g208(.A(G176gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT88), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT88), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n419_), .B(new_n420_), .C1(G183gat), .C2(G190gat), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n412_), .A2(new_n415_), .A3(new_n416_), .A4(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(G183gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(KEYINPUT25), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT26), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(G190gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427_));
  OAI22_X1  g226(.A1(KEYINPUT86), .A2(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT85), .B1(new_n429_), .B2(G183gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n423_), .A3(KEYINPUT25), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(KEYINPUT86), .A3(G183gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G190gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT26), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n425_), .A2(G190gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT87), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n428_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n406_), .A2(new_n410_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(KEYINPUT24), .A3(new_n416_), .ZN(new_n441_));
  OR3_X1    g240(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(new_n419_), .A3(new_n420_), .A4(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n422_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT20), .B1(new_n405_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n390_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G197gat), .B(G204gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n394_), .B1(new_n447_), .B2(new_n388_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n402_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n421_), .A2(new_n416_), .A3(new_n411_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT96), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n436_), .A2(new_n437_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n452_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT95), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n429_), .A2(G183gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n456_), .B1(new_n424_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n429_), .A2(G183gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n423_), .A2(KEYINPUT25), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(KEYINPUT95), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n443_), .B1(new_n455_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n451_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT26), .B(G190gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n452_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n435_), .A2(KEYINPUT26), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT96), .B1(new_n426_), .B2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n459_), .A2(new_n460_), .A3(KEYINPUT95), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT95), .B1(new_n459_), .B2(new_n460_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n467_), .B(new_n469_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n472_));
  AND4_X1   g271(.A1(new_n419_), .A2(new_n441_), .A3(new_n420_), .A4(new_n442_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT97), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n450_), .B1(new_n465_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n382_), .B1(new_n445_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT18), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n451_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n472_), .A2(new_n473_), .A3(new_n464_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n475_), .A2(new_n450_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n382_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n449_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n395_), .A2(KEYINPUT94), .A3(new_n402_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n444_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n485_), .A2(KEYINPUT20), .A3(new_n486_), .A4(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n477_), .A2(new_n482_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n482_), .B1(new_n477_), .B2(new_n491_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n380_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT102), .ZN(new_n495_));
  INV_X1    g294(.A(new_n491_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n488_), .A2(new_n489_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n434_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n500_), .A2(new_n459_), .B1(new_n436_), .B2(KEYINPUT87), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n499_), .B(new_n501_), .C1(KEYINPUT87), .C2(new_n466_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n412_), .A2(new_n415_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n421_), .A2(new_n416_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n502_), .A2(new_n473_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n497_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n484_), .A2(new_n483_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n464_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n449_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n486_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n481_), .B1(new_n496_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n477_), .A2(new_n482_), .A3(new_n491_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT102), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n380_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n495_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n490_), .A2(KEYINPUT20), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n463_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n382_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n506_), .A2(new_n509_), .A3(new_n486_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n481_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT27), .A3(new_n512_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526_));
  INV_X1    g325(.A(G155gat), .ZN(new_n527_));
  INV_X1    g326(.A(G162gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT90), .B1(G155gat), .B2(G162gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G155gat), .A2(G162gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT3), .ZN(new_n536_));
  INV_X1    g335(.A(G141gat), .ZN(new_n537_));
  INV_X1    g336(.A(G148gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n532_), .B1(new_n535_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n531_), .A2(KEYINPUT1), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT1), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(G155gat), .A3(G162gat), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n529_), .A2(new_n544_), .A3(new_n546_), .A4(new_n530_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G141gat), .B(G148gat), .Z(new_n548_));
  AND2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n525_), .B1(new_n543_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n532_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G141gat), .A2(G148gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT2), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n534_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n533_), .A2(KEYINPUT91), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n551_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n547_), .A2(new_n548_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(KEYINPUT92), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n550_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n524_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  AOI211_X1 g363(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n550_), .C2(new_n561_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G22gat), .B(G50gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n564_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n543_), .A2(new_n549_), .A3(new_n525_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT92), .B1(new_n559_), .B2(new_n560_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n563_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT28), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n562_), .A2(new_n524_), .A3(new_n563_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n566_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G78gat), .B(G106gat), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n541_), .A2(new_n540_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(new_n555_), .A3(new_n539_), .A4(new_n556_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n577_), .A2(new_n551_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n449_), .B1(new_n578_), .B2(new_n563_), .ZN(new_n579_));
  AND2_X1   g378(.A1(G228gat), .A2(G233gat), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n403_), .A2(new_n404_), .A3(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n550_), .A2(KEYINPUT29), .A3(new_n561_), .ZN(new_n582_));
  AOI221_X4 g381(.A(new_n575_), .B1(new_n579_), .B2(new_n580_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n575_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n580_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OAI22_X1  g386(.A1(new_n568_), .A2(new_n574_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n575_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n572_), .A2(new_n573_), .A3(new_n566_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n567_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n585_), .A2(new_n586_), .A3(new_n584_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .A4(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n516_), .A2(new_n523_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G71gat), .B(G99gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(G43gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n444_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G127gat), .B(G134gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G113gat), .B(G120gat), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(KEYINPUT89), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT89), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n602_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n600_), .B(new_n608_), .Z(new_n609_));
  NAND2_X1  g408(.A1(G227gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n351_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT30), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT31), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n609_), .B(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n550_), .A2(new_n561_), .A3(new_n608_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n603_), .A2(new_n604_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n578_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G225gat), .A2(G233gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G1gat), .B(G29gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G57gat), .B(G85gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n615_), .A2(KEYINPUT4), .A3(new_n617_), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT98), .B(KEYINPUT4), .Z(new_n626_));
  NAND4_X1  g425(.A1(new_n550_), .A2(new_n561_), .A3(new_n608_), .A4(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n618_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n619_), .B(new_n624_), .C1(new_n625_), .C2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT101), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n619_), .B1(new_n625_), .B2(new_n629_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n624_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n615_), .A2(new_n617_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT4), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n628_), .B(new_n627_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n619_), .A4(new_n624_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n631_), .A2(new_n634_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n614_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n597_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n514_), .B1(new_n513_), .B2(new_n380_), .ZN(new_n643_));
  AOI211_X1 g442(.A(KEYINPUT102), .B(KEYINPUT27), .C1(new_n511_), .C2(new_n512_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(new_n523_), .A3(new_n595_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT103), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n595_), .A2(new_n523_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n631_), .A2(new_n634_), .A3(new_n639_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n516_), .A3(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n492_), .A2(new_n493_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n630_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT33), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n630_), .A2(new_n654_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n635_), .A2(new_n628_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n659_), .B(new_n627_), .C1(new_n636_), .C2(new_n619_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n633_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n653_), .A2(new_n656_), .A3(new_n658_), .A4(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n496_), .A2(new_n510_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT32), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(new_n481_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n521_), .A2(KEYINPUT32), .A3(new_n482_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n649_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n662_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n596_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n647_), .A2(new_n652_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n614_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n642_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT83), .ZN(new_n673_));
  NAND2_X1  g472(.A1(G229gat), .A2(G233gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT82), .B1(new_n360_), .B2(new_n301_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT82), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n299_), .B(new_n676_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n355_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n357_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n356_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n350_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n301_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT81), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT81), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n682_), .A2(new_n301_), .A3(new_n686_), .A4(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n674_), .B1(new_n678_), .B2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n300_), .B(new_n303_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n688_), .A2(new_n674_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n673_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT84), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(new_n690_), .A3(new_n674_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n675_), .A2(new_n677_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n694_), .B(KEYINPUT83), .C1(new_n695_), .C2(new_n674_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(G113gat), .B(G141gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(G169gat), .B(G197gat), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n697_), .B(new_n698_), .Z(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n692_), .A2(new_n693_), .A3(new_n696_), .A4(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n694_), .B(new_n699_), .C1(new_n695_), .C2(new_n674_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n692_), .A2(new_n696_), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT84), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n672_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n379_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT80), .B1(new_n286_), .B2(new_n378_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n202_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n710_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n712_), .A2(KEYINPUT104), .A3(new_n708_), .A4(new_n379_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n640_), .A2(G1gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(KEYINPUT38), .A3(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n324_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT105), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n719_), .B(new_n324_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n672_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n284_), .A2(new_n707_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n375_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G1gat), .B1(new_n724_), .B2(new_n640_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n711_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT38), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n716_), .A2(new_n725_), .A3(new_n728_), .ZN(G1324gat));
  NAND2_X1  g528(.A1(new_n516_), .A2(new_n523_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(G8gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n711_), .A2(new_n713_), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G8gat), .B1(new_n724_), .B2(new_n731_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT39), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n734_), .A2(new_n735_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n733_), .A2(new_n736_), .A3(new_n737_), .A4(new_n739_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1325gat));
  NOR2_X1   g542(.A1(new_n671_), .A2(G15gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n714_), .A2(KEYINPUT107), .A3(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n711_), .A2(new_n713_), .A3(new_n744_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G15gat), .B1(new_n724_), .B2(new_n671_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT41), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n748_), .A3(new_n750_), .ZN(G1326gat));
  NAND3_X1  g550(.A1(new_n714_), .A2(new_n352_), .A3(new_n595_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G22gat), .B1(new_n724_), .B2(new_n596_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1327gat));
  NAND2_X1  g555(.A1(new_n721_), .A2(new_n374_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(new_n284_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n708_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G29gat), .B1(new_n760_), .B2(new_n649_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n346_), .A2(new_n377_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT43), .B1(new_n672_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n380_), .B1(new_n663_), .B2(new_n482_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n766_), .A2(new_n522_), .B1(new_n594_), .B2(new_n588_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n640_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n768_), .A2(KEYINPUT103), .B1(new_n668_), .B2(new_n596_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n614_), .B1(new_n769_), .B2(new_n652_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n765_), .B(new_n762_), .C1(new_n770_), .C2(new_n642_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n764_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n723_), .A2(new_n374_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT44), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n776_), .B(new_n773_), .C1(new_n764_), .C2(new_n771_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n649_), .A2(G29gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n761_), .B1(new_n778_), .B2(new_n779_), .ZN(G1328gat));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n781_));
  INV_X1    g580(.A(G36gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n778_), .B2(new_n730_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n731_), .A2(G36gat), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OR3_X1    g585(.A1(new_n759_), .A2(new_n784_), .A3(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n759_), .B2(new_n786_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n781_), .B1(new_n783_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n789_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n775_), .A2(new_n777_), .A3(new_n731_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n791_), .B(KEYINPUT46), .C1(new_n792_), .C2(new_n782_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(G1329gat));
  AOI21_X1  g593(.A(G43gat), .B1(new_n760_), .B2(new_n614_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n614_), .A2(G43gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n778_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n798_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n795_), .B(new_n800_), .C1(new_n778_), .C2(new_n796_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1330gat));
  NAND2_X1  g601(.A1(new_n772_), .A2(new_n774_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n776_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n772_), .A2(KEYINPUT44), .A3(new_n774_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n595_), .A3(new_n805_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT111), .B1(new_n806_), .B2(G50gat), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n596_), .A2(G50gat), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT112), .Z(new_n810_));
  OAI22_X1  g609(.A1(new_n807_), .A2(new_n808_), .B1(new_n759_), .B2(new_n810_), .ZN(G1331gat));
  NAND2_X1  g610(.A1(new_n378_), .A2(new_n284_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(KEYINPUT113), .Z(new_n813_));
  NOR2_X1   g612(.A1(new_n672_), .A2(new_n706_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(KEYINPUT114), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n812_), .B(KEYINPUT113), .ZN(new_n817_));
  INV_X1    g616(.A(new_n814_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(G57gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n649_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n282_), .A2(new_n283_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(KEYINPUT71), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n284_), .A2(new_n285_), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n374_), .A4(new_n706_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n722_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G57gat), .B1(new_n827_), .B2(new_n640_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n822_), .A2(new_n828_), .ZN(G1332gat));
  INV_X1    g628(.A(G64gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n820_), .A2(new_n830_), .A3(new_n730_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G64gat), .B1(new_n827_), .B2(new_n731_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n832_), .A2(KEYINPUT48), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(KEYINPUT48), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n831_), .B1(new_n833_), .B2(new_n834_), .ZN(G1333gat));
  OAI21_X1  g634(.A(G71gat), .B1(new_n827_), .B2(new_n671_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT116), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n671_), .A2(G71gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n815_), .A2(new_n819_), .A3(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(G71gat), .B(new_n838_), .C1(new_n827_), .C2(new_n671_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT117), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n840_), .A2(new_n842_), .A3(new_n846_), .A4(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1334gat));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n849_));
  OAI21_X1  g648(.A(G78gat), .B1(new_n827_), .B2(new_n596_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT118), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(KEYINPUT118), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n849_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n850_), .A2(KEYINPUT118), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(KEYINPUT50), .A3(new_n851_), .ZN(new_n856_));
  INV_X1    g655(.A(G78gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n820_), .A2(new_n857_), .A3(new_n595_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(new_n856_), .A3(new_n858_), .ZN(G1335gat));
  NOR2_X1   g658(.A1(new_n375_), .A2(new_n706_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n284_), .A2(KEYINPUT119), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT119), .B1(new_n284_), .B2(new_n860_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n764_), .B2(new_n771_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G85gat), .B1(new_n865_), .B2(new_n640_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n818_), .A2(new_n286_), .A3(new_n757_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n214_), .A3(new_n649_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1336gat));
  OAI21_X1  g668(.A(G92gat), .B1(new_n865_), .B2(new_n731_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n867_), .A2(new_n215_), .A3(new_n730_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1337gat));
  NAND3_X1  g671(.A1(new_n867_), .A2(new_n224_), .A3(new_n614_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n865_), .A2(new_n671_), .ZN(new_n874_));
  INV_X1    g673(.A(G99gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n876_), .B(new_n878_), .ZN(G1338gat));
  NAND3_X1  g678(.A1(new_n867_), .A2(new_n225_), .A3(new_n595_), .ZN(new_n880_));
  AOI211_X1 g679(.A(KEYINPUT52), .B(new_n225_), .C1(new_n864_), .C2(new_n595_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n882_));
  INV_X1    g681(.A(new_n863_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n772_), .A2(new_n595_), .A3(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n884_), .B2(G106gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n880_), .B1(new_n881_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT53), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n888_), .B(new_n880_), .C1(new_n881_), .C2(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1339gat));
  OAI21_X1  g689(.A(KEYINPUT55), .B1(new_n256_), .B2(KEYINPUT121), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT55), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n261_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n244_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n247_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n891_), .A2(new_n894_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n270_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n897_), .A2(KEYINPUT56), .A3(new_n270_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n674_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n688_), .A2(new_n690_), .A3(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n904_), .B(new_n700_), .C1(new_n695_), .C2(new_n903_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n702_), .A2(new_n905_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n278_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n902_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n902_), .A2(KEYINPUT58), .A3(new_n907_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n762_), .A3(new_n911_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n703_), .A2(new_n705_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n901_), .ZN(new_n914_));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n897_), .B2(new_n270_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n280_), .A2(new_n906_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n721_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT57), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n912_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n918_), .A2(KEYINPUT57), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n374_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n282_), .A2(new_n283_), .A3(new_n707_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(new_n378_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n282_), .A2(new_n283_), .A3(new_n707_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n346_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n926_), .A2(new_n927_), .A3(KEYINPUT54), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n925_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n922_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n597_), .A2(new_n640_), .A3(new_n671_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT122), .B1(new_n918_), .B2(KEYINPUT57), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n902_), .A2(new_n913_), .B1(new_n280_), .B2(new_n906_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n936_), .B(new_n937_), .C1(new_n938_), .C2(new_n721_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n935_), .A2(new_n939_), .A3(new_n912_), .A4(new_n919_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n929_), .B1(new_n940_), .B2(new_n374_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n933_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n934_), .B1(new_n943_), .B2(new_n932_), .ZN(new_n944_));
  OAI21_X1  g743(.A(G113gat), .B1(new_n944_), .B2(new_n707_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n943_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n707_), .A2(G113gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n945_), .B1(new_n946_), .B2(new_n947_), .ZN(G1340gat));
  OAI21_X1  g747(.A(G120gat), .B1(new_n944_), .B2(new_n286_), .ZN(new_n949_));
  INV_X1    g748(.A(G120gat), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n950_), .B1(new_n823_), .B2(KEYINPUT60), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n951_), .B1(KEYINPUT60), .B2(new_n950_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n949_), .B1(new_n946_), .B2(new_n952_), .ZN(G1341gat));
  OAI21_X1  g752(.A(G127gat), .B1(new_n944_), .B2(new_n374_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n374_), .A2(G127gat), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n946_), .B2(new_n955_), .ZN(G1342gat));
  OAI21_X1  g755(.A(G134gat), .B1(new_n944_), .B2(new_n763_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n721_), .ZN(new_n958_));
  OR2_X1    g757(.A1(new_n958_), .A2(G134gat), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n946_), .B2(new_n959_), .ZN(G1343gat));
  NOR2_X1   g759(.A1(new_n614_), .A2(new_n596_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n941_), .A2(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n730_), .A2(new_n640_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n963_), .A2(new_n706_), .A3(new_n964_), .ZN(new_n965_));
  XOR2_X1   g764(.A(KEYINPUT123), .B(G141gat), .Z(new_n966_));
  XNOR2_X1  g765(.A(new_n965_), .B(new_n966_), .ZN(G1344gat));
  NOR2_X1   g766(.A1(new_n824_), .A2(new_n825_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n963_), .A2(new_n968_), .A3(new_n964_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g769(.A1(new_n963_), .A2(new_n375_), .A3(new_n964_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(KEYINPUT61), .B(G155gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n971_), .B(new_n972_), .ZN(G1346gat));
  INV_X1    g772(.A(new_n941_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n958_), .A2(G162gat), .ZN(new_n975_));
  NAND4_X1  g774(.A1(new_n974_), .A2(new_n961_), .A3(new_n964_), .A4(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(new_n964_), .ZN(new_n977_));
  NOR4_X1   g776(.A1(new_n941_), .A2(new_n763_), .A3(new_n962_), .A4(new_n977_), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n976_), .B1(new_n978_), .B2(new_n528_), .ZN(new_n979_));
  INV_X1    g778(.A(KEYINPUT124), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(new_n981_));
  OAI211_X1 g780(.A(new_n976_), .B(KEYINPUT124), .C1(new_n978_), .C2(new_n528_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(G1347gat));
  NOR2_X1   g782(.A1(new_n731_), .A2(new_n649_), .ZN(new_n984_));
  INV_X1    g783(.A(new_n984_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n985_), .A2(new_n671_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(new_n596_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n987_), .B1(new_n922_), .B2(new_n930_), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n406_), .B1(new_n988_), .B2(new_n706_), .ZN(new_n989_));
  OR2_X1    g788(.A1(new_n989_), .A2(KEYINPUT62), .ZN(new_n990_));
  NAND3_X1  g789(.A1(new_n988_), .A2(new_n413_), .A3(new_n706_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n989_), .A2(KEYINPUT62), .ZN(new_n992_));
  NAND3_X1  g791(.A1(new_n990_), .A2(new_n991_), .A3(new_n992_), .ZN(G1348gat));
  AOI21_X1  g792(.A(G176gat), .B1(new_n988_), .B2(new_n284_), .ZN(new_n994_));
  NOR2_X1   g793(.A1(new_n941_), .A2(new_n595_), .ZN(new_n995_));
  INV_X1    g794(.A(new_n986_), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n996_), .A2(new_n410_), .A3(new_n286_), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n994_), .B1(new_n995_), .B2(new_n997_), .ZN(G1349gat));
  NOR4_X1   g797(.A1(new_n941_), .A2(new_n374_), .A3(new_n595_), .A4(new_n996_), .ZN(new_n999_));
  OR2_X1    g798(.A1(new_n999_), .A2(KEYINPUT125), .ZN(new_n1000_));
  AOI21_X1  g799(.A(G183gat), .B1(new_n999_), .B2(KEYINPUT125), .ZN(new_n1001_));
  NOR2_X1   g800(.A1(new_n374_), .A2(new_n462_), .ZN(new_n1002_));
  AOI22_X1  g801(.A1(new_n1000_), .A2(new_n1001_), .B1(new_n988_), .B2(new_n1002_), .ZN(G1350gat));
  AND2_X1   g802(.A1(new_n721_), .A2(new_n455_), .ZN(new_n1004_));
  AND2_X1   g803(.A1(new_n988_), .A2(new_n1004_), .ZN(new_n1005_));
  AOI21_X1  g804(.A(new_n435_), .B1(new_n988_), .B2(new_n762_), .ZN(new_n1006_));
  NOR2_X1   g805(.A1(new_n1005_), .A2(new_n1006_), .ZN(new_n1007_));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1008_));
  NAND2_X1  g807(.A1(new_n1007_), .A2(new_n1008_), .ZN(new_n1009_));
  OAI21_X1  g808(.A(KEYINPUT126), .B1(new_n1005_), .B2(new_n1006_), .ZN(new_n1010_));
  NAND2_X1  g809(.A1(new_n1009_), .A2(new_n1010_), .ZN(G1351gat));
  NAND3_X1  g810(.A1(new_n963_), .A2(new_n706_), .A3(new_n984_), .ZN(new_n1012_));
  XNOR2_X1  g811(.A(new_n1012_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g812(.A1(new_n963_), .A2(new_n968_), .A3(new_n984_), .ZN(new_n1014_));
  XNOR2_X1  g813(.A(new_n1014_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g814(.A(new_n374_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1016_));
  NOR2_X1   g815(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1017_));
  NAND2_X1  g816(.A1(new_n1017_), .A2(KEYINPUT127), .ZN(new_n1018_));
  AND4_X1   g817(.A1(new_n963_), .A2(new_n984_), .A3(new_n1016_), .A4(new_n1018_), .ZN(new_n1019_));
  NAND2_X1  g818(.A1(new_n974_), .A2(new_n961_), .ZN(new_n1020_));
  NOR2_X1   g819(.A1(new_n1020_), .A2(new_n985_), .ZN(new_n1021_));
  NAND2_X1  g820(.A1(new_n1021_), .A2(new_n1016_), .ZN(new_n1022_));
  XNOR2_X1  g821(.A(new_n1017_), .B(KEYINPUT127), .ZN(new_n1023_));
  AOI21_X1  g822(.A(new_n1019_), .B1(new_n1022_), .B2(new_n1023_), .ZN(G1354gat));
  NAND3_X1  g823(.A1(new_n1021_), .A2(new_n397_), .A3(new_n721_), .ZN(new_n1025_));
  NOR3_X1   g824(.A1(new_n1020_), .A2(new_n763_), .A3(new_n985_), .ZN(new_n1026_));
  OAI21_X1  g825(.A(new_n1025_), .B1(new_n397_), .B2(new_n1026_), .ZN(G1355gat));
endmodule


