//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(KEYINPUT9), .A3(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n204_), .A2(new_n209_), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  OAI22_X1  g016(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .A4(new_n203_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n207_), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n218_), .B(new_n222_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT66), .B1(new_n213_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n210_), .A2(new_n228_), .A3(new_n211_), .ZN(new_n229_));
  AND4_X1   g028(.A1(new_n217_), .A2(new_n225_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n227_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n217_), .B1(new_n231_), .B2(new_n225_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n216_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G71gat), .B(G78gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G57gat), .A2(G64gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G57gat), .A2(G64gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT67), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G57gat), .ZN(new_n240_));
  INV_X1    g039(.A(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n236_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n235_), .B1(new_n245_), .B2(KEYINPUT11), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n239_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(KEYINPUT11), .A3(new_n235_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n233_), .A2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n209_), .A2(new_n218_), .A3(new_n222_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n229_), .A2(new_n227_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT8), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n231_), .A2(new_n217_), .A3(new_n225_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AOI211_X1 g056(.A(new_n248_), .B(new_n234_), .C1(new_n239_), .C2(new_n244_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n246_), .A2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n257_), .A2(new_n259_), .A3(new_n216_), .A4(new_n249_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n252_), .A2(new_n260_), .A3(KEYINPUT12), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n233_), .A2(new_n251_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G230gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT64), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n252_), .A2(new_n260_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n266_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G176gat), .B(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G148gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT69), .B(G120gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n267_), .A2(new_n270_), .A3(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n281_), .A2(KEYINPUT13), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(KEYINPUT13), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT70), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(KEYINPUT70), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT84), .ZN(new_n289_));
  INV_X1    g088(.A(G50gat), .ZN(new_n290_));
  OR2_X1    g089(.A1(G29gat), .A2(G36gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G29gat), .A2(G36gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n295_), .A2(G43gat), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G43gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G29gat), .B(G36gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT71), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n300_), .B2(new_n294_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n290_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(G43gat), .B1(new_n295_), .B2(new_n296_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n298_), .A3(new_n294_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(G50gat), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT77), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G15gat), .B(G22gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n312_), .B(KEYINPUT14), .C1(new_n307_), .C2(new_n308_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G1gat), .B(G8gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n306_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT15), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n297_), .A2(new_n301_), .A3(new_n290_), .ZN(new_n319_));
  AOI21_X1  g118(.A(G50gat), .B1(new_n303_), .B2(new_n304_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n302_), .A2(KEYINPUT15), .A3(new_n305_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n316_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n317_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G229gat), .A2(G233gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT83), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n306_), .B(new_n324_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n330_), .A2(new_n326_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G141gat), .ZN(new_n333_));
  INV_X1    g132(.A(G169gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G197gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n289_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n329_), .A2(new_n331_), .A3(KEYINPUT84), .A4(new_n339_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n338_), .A2(new_n340_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n288_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G71gat), .B(G99gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT23), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G183gat), .A3(G190gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT88), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT88), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n349_), .B2(KEYINPUT23), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n348_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT86), .ZN(new_n360_));
  INV_X1    g159(.A(G176gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G169gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OAI221_X1 g162(.A(KEYINPUT89), .B1(G183gat), .B2(G190gat), .C1(new_n353_), .C2(new_n355_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n358_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT30), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n360_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n350_), .A2(new_n352_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT24), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n334_), .A3(new_n361_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(KEYINPUT87), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n376_));
  INV_X1    g175(.A(G190gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(KEYINPUT26), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT25), .B(G183gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT26), .B(G190gat), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n378_), .B(new_n379_), .C1(new_n380_), .C2(new_n376_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n368_), .A2(new_n372_), .A3(new_n375_), .A4(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n365_), .A2(new_n366_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n366_), .B1(new_n365_), .B2(new_n382_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n347_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n365_), .A2(new_n382_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT30), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n365_), .A2(new_n366_), .A3(new_n382_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT31), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G113gat), .B(G120gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(KEYINPUT90), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n390_), .B(new_n391_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(KEYINPUT90), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G15gat), .B(G43gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n385_), .A2(new_n389_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n385_), .B2(new_n389_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n346_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n385_), .A2(new_n389_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n397_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n385_), .A2(new_n389_), .A3(new_n397_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n345_), .A3(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT98), .ZN(new_n408_));
  OR2_X1    g207(.A1(G155gat), .A2(G162gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT2), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n409_), .B(new_n410_), .C1(new_n413_), .C2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n411_), .B(KEYINPUT91), .ZN(new_n418_));
  AND3_X1   g217(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n409_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n421_), .A3(new_n414_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT29), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G228gat), .A2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G211gat), .B(G218gat), .Z(new_n427_));
  INV_X1    g226(.A(KEYINPUT94), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n336_), .B2(G204gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n336_), .A2(G204gat), .ZN(new_n430_));
  INV_X1    g229(.A(G204gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(KEYINPUT94), .A3(G197gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n427_), .B1(new_n433_), .B2(KEYINPUT21), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n435_), .A2(KEYINPUT21), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n431_), .A2(G197gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(KEYINPUT21), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n430_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n430_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n427_), .A2(KEYINPUT21), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n426_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n424_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT96), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n424_), .A2(new_n444_), .A3(KEYINPUT96), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(new_n443_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT97), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n442_), .B1(new_n434_), .B2(new_n439_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT97), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n454_), .A3(new_n424_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n426_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n408_), .B1(new_n449_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n417_), .A2(new_n458_), .A3(new_n422_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT92), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G22gat), .B(G50gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n461_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(new_n417_), .A3(new_n458_), .A4(new_n422_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n464_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n407_), .B1(new_n457_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n407_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n447_), .A2(new_n448_), .B1(new_n455_), .B2(new_n426_), .ZN(new_n472_));
  OAI221_X1 g271(.A(new_n471_), .B1(new_n467_), .B2(new_n468_), .C1(new_n472_), .C2(new_n408_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n408_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n475_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n470_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n406_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n400_), .A2(new_n405_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n470_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n477_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n371_), .A2(new_n367_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT99), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT99), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n371_), .A2(new_n487_), .A3(new_n367_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n359_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n380_), .A2(new_n379_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n489_), .B(new_n490_), .C1(new_n353_), .C2(new_n355_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n369_), .B1(G183gat), .B2(G190gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n363_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n450_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n365_), .A2(new_n382_), .A3(new_n453_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G226gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT19), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT20), .A4(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n494_), .A2(new_n450_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n453_), .B1(new_n365_), .B2(new_n382_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n499_), .B1(new_n503_), .B2(new_n498_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n499_), .B(new_n509_), .C1(new_n503_), .C2(new_n498_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT104), .B(KEYINPUT27), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(new_n504_), .B2(new_n510_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n495_), .A2(KEYINPUT20), .A3(new_n496_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(new_n498_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n494_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT102), .B1(new_n520_), .B2(new_n502_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT102), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n453_), .B(new_n451_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n522_), .B(KEYINPUT20), .C1(new_n523_), .C2(new_n494_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n501_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n519_), .B1(new_n526_), .B2(new_n498_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n509_), .B(KEYINPUT103), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n517_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G225gat), .A2(G233gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n395_), .A2(new_n423_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n417_), .A2(new_n394_), .A3(new_n422_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT4), .B1(new_n395_), .B2(new_n423_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n531_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G1gat), .B(G29gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G85gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT0), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n240_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n533_), .A2(new_n530_), .A3(new_n534_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n537_), .B2(new_n542_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n515_), .A2(new_n529_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n484_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n544_), .A2(new_n545_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n510_), .A2(KEYINPUT32), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n504_), .A2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n550_), .B(new_n552_), .C1(new_n527_), .C2(new_n551_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT33), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT101), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n543_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n541_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n530_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n533_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n556_), .A2(new_n511_), .A3(new_n512_), .A4(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n476_), .A2(new_n478_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n406_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n549_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n342_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n321_), .A2(new_n322_), .A3(new_n233_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT34), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(KEYINPUT35), .A3(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(KEYINPUT35), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT72), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n306_), .A2(new_n257_), .A3(new_n216_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n573_), .A2(KEYINPUT72), .ZN(new_n576_));
  AND4_X1   g375(.A1(new_n567_), .A2(new_n574_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n567_), .A2(new_n574_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n571_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT74), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G134gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G162gat), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(KEYINPUT36), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n578_), .A2(new_n588_), .A3(new_n582_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n587_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT76), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n600_), .B2(KEYINPUT37), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT76), .B(new_n602_), .C1(new_n591_), .C2(new_n599_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n597_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n595_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(KEYINPUT37), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT76), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n600_), .A2(new_n598_), .A3(KEYINPUT37), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n605_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n604_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT78), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n316_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n251_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n615_), .A2(KEYINPUT79), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(KEYINPUT79), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT81), .ZN(new_n619_));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT17), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n616_), .A2(new_n617_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n624_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n615_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT82), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT82), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n615_), .A2(new_n625_), .A3(new_n630_), .A4(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n626_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n611_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n566_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n307_), .A3(new_n550_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT38), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n634_), .A2(new_n597_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n566_), .A2(new_n550_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G1gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(G1324gat));
  NAND2_X1  g441(.A1(new_n515_), .A2(new_n529_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(new_n308_), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n566_), .A2(new_n643_), .A3(new_n639_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(G8gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n645_), .B2(G8gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n644_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n636_), .A2(new_n653_), .A3(new_n480_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n566_), .A2(new_n480_), .A3(new_n639_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT41), .B1(new_n655_), .B2(G15gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT105), .ZN(G1326gat));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n563_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n636_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n566_), .A2(new_n662_), .A3(new_n639_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(G22gat), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n665_), .B1(new_n664_), .B2(G22gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT107), .ZN(G1327gat));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n607_), .A2(new_n605_), .A3(new_n608_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n597_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n549_), .A2(new_n564_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n675_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n406_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n553_), .B2(new_n561_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n547_), .B1(new_n479_), .B2(new_n483_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT109), .B(new_n677_), .C1(new_n610_), .C2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n674_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n676_), .A2(new_n682_), .A3(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n342_), .A3(new_n634_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n687_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n550_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G29gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n633_), .A2(new_n605_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n342_), .A2(new_n565_), .A3(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n546_), .A2(G29gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(new_n643_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n693_), .A2(G36gat), .A3(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT45), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n688_), .A2(new_n643_), .A3(new_n689_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n700_), .A3(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  NAND3_X1  g504(.A1(new_n688_), .A2(new_n480_), .A3(new_n689_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G43gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n693_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n298_), .A3(new_n480_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(KEYINPUT47), .A3(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1330gat));
  NAND3_X1  g513(.A1(new_n708_), .A2(new_n290_), .A3(new_n662_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n688_), .A2(new_n662_), .A3(new_n689_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(new_n290_), .ZN(G1331gat));
  INV_X1    g516(.A(new_n341_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n287_), .A2(new_n718_), .A3(new_n681_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n639_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n240_), .A3(new_n546_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n719_), .A2(new_n635_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n722_), .A2(KEYINPUT110), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(KEYINPUT110), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n550_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n721_), .B1(new_n725_), .B2(new_n240_), .ZN(G1332gat));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n241_), .A3(new_n643_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728_));
  INV_X1    g527(.A(new_n720_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n643_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n730_), .B2(G64gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT48), .B(new_n241_), .C1(new_n729_), .C2(new_n643_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT111), .Z(G1333gat));
  INV_X1    g533(.A(G71gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n722_), .A2(new_n735_), .A3(new_n480_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G71gat), .B1(new_n720_), .B2(new_n406_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n737_), .A2(new_n738_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1334gat));
  OAI21_X1  g540(.A(G78gat), .B1(new_n720_), .B2(new_n563_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT50), .ZN(new_n743_));
  INV_X1    g542(.A(G78gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n722_), .A2(new_n744_), .A3(new_n662_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1335gat));
  AND2_X1   g545(.A1(new_n719_), .A2(new_n692_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n550_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n685_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n287_), .A2(new_n718_), .A3(new_n633_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n550_), .A2(G85gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT113), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n748_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT114), .ZN(G1336gat));
  INV_X1    g555(.A(G92gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n747_), .A2(new_n757_), .A3(new_n643_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n749_), .A2(new_n696_), .A3(new_n751_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n757_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT115), .ZN(G1337gat));
  NAND3_X1  g560(.A1(new_n747_), .A2(new_n202_), .A3(new_n480_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n749_), .A2(new_n406_), .A3(new_n751_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n221_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n764_), .B(new_n765_), .Z(G1338gat));
  NAND3_X1  g565(.A1(new_n685_), .A2(new_n662_), .A3(new_n750_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT117), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n685_), .A2(new_n769_), .A3(new_n662_), .A4(new_n750_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(G106gat), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT52), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n768_), .A2(new_n773_), .A3(G106gat), .A4(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n747_), .A2(new_n203_), .A3(new_n662_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n779_), .A3(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  OAI211_X1 g580(.A(new_n633_), .B(new_n341_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n610_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT120), .Z(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n784_), .A2(new_n610_), .A3(new_n787_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n267_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n264_), .A2(KEYINPUT55), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n269_), .A2(KEYINPUT121), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n264_), .A2(KEYINPUT55), .A3(new_n795_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT122), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT122), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n793_), .A2(new_n797_), .A3(new_n801_), .A4(new_n798_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n278_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n278_), .A4(new_n802_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT123), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n280_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n341_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT123), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n803_), .A2(new_n810_), .A3(new_n804_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n330_), .A2(new_n327_), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n339_), .B(new_n813_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n281_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n597_), .B1(new_n812_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT57), .B1(new_n817_), .B2(KEYINPUT124), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n805_), .A2(new_n806_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(new_n280_), .A3(new_n815_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n819_), .A2(KEYINPUT58), .A3(new_n280_), .A4(new_n815_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n611_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n811_), .A2(new_n809_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n827_), .A2(new_n807_), .B1(new_n281_), .B2(new_n815_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n825_), .B(new_n826_), .C1(new_n828_), .C2(new_n597_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n818_), .A2(new_n824_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n791_), .B1(new_n830_), .B2(new_n634_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n643_), .A2(new_n546_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n831_), .A2(new_n483_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834_), .B2(new_n718_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n830_), .A2(new_n634_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n791_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT125), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT59), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n476_), .A2(new_n478_), .B1(new_n405_), .B2(new_n400_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n841_), .A3(new_n832_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n831_), .B2(KEYINPUT125), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n834_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n341_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n835_), .B1(new_n847_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n287_), .B2(KEYINPUT60), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(KEYINPUT60), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(KEYINPUT126), .B2(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n834_), .B(new_n852_), .C1(KEYINPUT126), .C2(new_n850_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n287_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n849_), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n834_), .B2(new_n633_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n634_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g657(.A(G134gat), .B1(new_n834_), .B2(new_n597_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n610_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g660(.A1(new_n831_), .A2(new_n479_), .A3(new_n833_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n718_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n288_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n633_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  AOI21_X1  g668(.A(G162gat), .B1(new_n862_), .B2(new_n597_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n611_), .A2(G162gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n862_), .B2(new_n871_), .ZN(G1347gat));
  AOI21_X1  g671(.A(new_n483_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n696_), .A2(new_n550_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n873_), .A2(new_n718_), .A3(new_n362_), .A4(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n874_), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n831_), .A2(new_n341_), .A3(new_n483_), .A4(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n334_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n877_), .B2(new_n334_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1348gat));
  NAND3_X1  g681(.A1(new_n873_), .A2(new_n288_), .A3(new_n874_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g683(.A1(new_n873_), .A2(new_n633_), .A3(new_n874_), .ZN(new_n885_));
  MUX2_X1   g684(.A(new_n379_), .B(G183gat), .S(new_n885_), .Z(G1350gat));
  NAND4_X1  g685(.A1(new_n873_), .A2(new_n380_), .A3(new_n597_), .A4(new_n874_), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n831_), .A2(new_n483_), .A3(new_n610_), .A4(new_n876_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n377_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n831_), .A2(new_n479_), .A3(new_n876_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n718_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n288_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n633_), .A3(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT127), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n896_), .B(new_n898_), .ZN(G1354gat));
  AOI21_X1  g698(.A(G218gat), .B1(new_n890_), .B2(new_n597_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n611_), .A2(G218gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n890_), .B2(new_n901_), .ZN(G1355gat));
endmodule


