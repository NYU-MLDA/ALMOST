//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(KEYINPUT9), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT10), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT10), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  AND3_X1   g012(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n217_));
  AND4_X1   g016(.A1(new_n207_), .A2(new_n213_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n205_), .A2(new_n206_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n211_), .A4(new_n208_), .ZN(new_n222_));
  OAI22_X1  g021(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n219_), .B1(new_n224_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n233_), .B(new_n219_), .C1(new_n224_), .C2(new_n230_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n218_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G43gat), .B(G50gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT71), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT70), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT71), .ZN(new_n240_));
  INV_X1    g039(.A(G29gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(G36gat), .ZN(new_n242_));
  INV_X1    g041(.A(G36gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(G29gat), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n238_), .B(new_n240_), .C1(new_n242_), .C2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n238_), .A2(new_n240_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n236_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n245_), .A2(new_n248_), .A3(new_n236_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT35), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n254_));
  NAND2_X1  g053(.A1(G232gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n235_), .A2(new_n252_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n213_), .A2(new_n207_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n216_), .A2(new_n229_), .A3(new_n223_), .A4(new_n222_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n233_), .B1(new_n259_), .B2(new_n219_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n234_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n258_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n250_), .A2(KEYINPUT15), .A3(new_n251_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT15), .ZN(new_n264_));
  INV_X1    g063(.A(new_n251_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(new_n249_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n263_), .A3(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n256_), .A2(new_n253_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n257_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n256_), .A2(new_n253_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n265_), .A2(new_n249_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n262_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n257_), .A2(KEYINPUT73), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n262_), .A2(new_n263_), .A3(new_n266_), .A4(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n267_), .A2(KEYINPUT72), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n268_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n270_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G190gat), .B(G218gat), .Z(new_n283_));
  XOR2_X1   g082(.A(G134gat), .B(G162gat), .Z(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n282_), .A2(KEYINPUT75), .A3(new_n285_), .A4(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n280_), .A2(new_n281_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n269_), .ZN(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n285_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT77), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT78), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT78), .ZN(new_n299_));
  INV_X1    g098(.A(new_n297_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n282_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n202_), .B1(new_n292_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n288_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n282_), .A2(new_n296_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n304_), .A2(new_n305_), .A3(KEYINPUT37), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT79), .B1(new_n303_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT79), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n294_), .A2(KEYINPUT78), .A3(new_n297_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n299_), .B1(new_n282_), .B2(new_n300_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n308_), .B1(new_n312_), .B2(new_n202_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G15gat), .B(G22gat), .ZN(new_n315_));
  INV_X1    g114(.A(G1gat), .ZN(new_n316_));
  INV_X1    g115(.A(G8gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT14), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G8gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G231gat), .A2(G233gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  XNOR2_X1  g122(.A(G57gat), .B(G64gat), .ZN(new_n324_));
  INV_X1    g123(.A(G71gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT65), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G71gat), .ZN(new_n328_));
  INV_X1    g127(.A(G78gat), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT11), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n327_), .A2(G71gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n325_), .A2(KEYINPUT65), .ZN(new_n335_));
  OAI21_X1  g134(.A(G78gat), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT11), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n324_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(KEYINPUT11), .A3(new_n337_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n324_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n323_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT17), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G155gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G211gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT16), .B(G183gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  OAI21_X1  g149(.A(new_n345_), .B1(new_n346_), .B2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n346_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n344_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n314_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT80), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G64gat), .B(G92gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G211gat), .B(G218gat), .Z(new_n363_));
  INV_X1    g162(.A(G197gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(KEYINPUT89), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(G204gat), .ZN(new_n366_));
  INV_X1    g165(.A(G204gat), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT90), .B(KEYINPUT21), .C1(new_n364_), .C2(new_n367_), .ZN(new_n368_));
  OR3_X1    g167(.A1(new_n363_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(G197gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT21), .ZN(new_n371_));
  OAI221_X1 g170(.A(new_n370_), .B1(new_n367_), .B2(new_n365_), .C1(new_n363_), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n364_), .A2(KEYINPUT89), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT90), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n363_), .B1(new_n374_), .B2(new_n371_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(new_n372_), .A3(new_n373_), .A4(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(G169gat), .B2(G176gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT25), .B(G183gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT26), .B(G190gat), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OR3_X1    g181(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384_));
  INV_X1    g183(.A(G183gat), .ZN(new_n385_));
  INV_X1    g184(.A(G190gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(KEYINPUT93), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT93), .ZN(new_n391_));
  AOI221_X4 g190(.A(new_n379_), .B1(new_n380_), .B2(new_n382_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n387_), .A2(new_n388_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(G183gat), .B2(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT22), .B(G169gat), .ZN(new_n398_));
  INV_X1    g197(.A(G176gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n377_), .B1(new_n392_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT19), .ZN(new_n405_));
  NAND2_X1  g204(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G169gat), .ZN(new_n407_));
  INV_X1    g206(.A(G169gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n409_), .A3(new_n399_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n397_), .A2(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n411_), .A2(KEYINPUT85), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(KEYINPUT85), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n394_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n378_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n397_), .A2(new_n415_), .ZN(new_n416_));
  OR3_X1    g215(.A1(new_n386_), .A2(KEYINPUT82), .A3(KEYINPUT26), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT26), .B1(new_n386_), .B2(KEYINPUT82), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n380_), .A3(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n383_), .A3(new_n393_), .A4(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n414_), .A2(new_n420_), .A3(new_n376_), .ZN(new_n421_));
  AND4_X1   g220(.A1(KEYINPUT20), .A2(new_n403_), .A3(new_n405_), .A4(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n376_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n379_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n382_), .A2(new_n380_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n376_), .A3(new_n401_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n405_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n362_), .B1(new_n422_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT95), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n403_), .A2(KEYINPUT20), .A3(new_n421_), .A4(new_n405_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n414_), .A2(new_n420_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n377_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n435_), .A2(KEYINPUT20), .A3(new_n429_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n361_), .B(new_n433_), .C1(new_n436_), .C2(new_n405_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n433_), .B1(new_n436_), .B2(new_n405_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(KEYINPUT95), .A3(new_n362_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G155gat), .A2(G162gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(G141gat), .A2(G148gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT3), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(KEYINPUT2), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G141gat), .A2(G148gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n447_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(new_n448_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n444_), .B1(new_n446_), .B2(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n442_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n444_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n445_), .B(new_n454_), .C1(new_n455_), .C2(KEYINPUT1), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G127gat), .B(G134gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G120gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n462_), .A2(KEYINPUT4), .A3(new_n464_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n464_), .A2(KEYINPUT4), .ZN(new_n469_));
  INV_X1    g268(.A(new_n466_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(new_n203_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT0), .B(G57gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT96), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(KEYINPUT96), .A3(KEYINPUT33), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n465_), .A2(new_n470_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n468_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n475_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n441_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n362_), .A2(KEYINPUT32), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n439_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT97), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n467_), .A2(new_n471_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n484_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n476_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n405_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n436_), .A2(new_n494_), .ZN(new_n495_));
  AND4_X1   g294(.A1(KEYINPUT20), .A2(new_n403_), .A3(new_n494_), .A4(new_n421_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT32), .B(new_n362_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n439_), .A2(KEYINPUT97), .A3(new_n487_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n490_), .A2(new_n493_), .A3(new_n497_), .A4(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n486_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G99gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G227gat), .A2(G233gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n414_), .A2(new_n504_), .A3(new_n420_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n463_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n434_), .A2(KEYINPUT30), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n461_), .A3(new_n505_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G15gat), .B(G43gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT31), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n513_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n503_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(new_n503_), .A3(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G78gat), .B(G106gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT91), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n376_), .B1(KEYINPUT29), .B2(new_n457_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(G228gat), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n457_), .A2(KEYINPUT29), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n531_), .A2(new_n377_), .A3(new_n529_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n524_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n377_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n529_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n525_), .A2(new_n529_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n523_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n538_), .A3(KEYINPUT92), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n536_), .A2(new_n537_), .A3(new_n540_), .A4(new_n523_), .ZN(new_n541_));
  INV_X1    g340(.A(G50gat), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n458_), .B2(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n457_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT28), .B(G22gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n544_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n458_), .A2(new_n543_), .A3(new_n542_), .ZN(new_n549_));
  OAI21_X1  g348(.A(G50gat), .B1(new_n457_), .B2(KEYINPUT29), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n548_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n547_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT87), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n539_), .B(new_n541_), .C1(new_n553_), .C2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n533_), .A2(new_n538_), .A3(new_n555_), .A4(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n500_), .A2(new_n521_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n519_), .A3(new_n518_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n516_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n515_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n503_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n557_), .B(new_n558_), .C1(new_n566_), .C2(new_n517_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT27), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n438_), .A2(new_n569_), .A3(new_n440_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n431_), .A2(KEYINPUT98), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT98), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n439_), .A2(new_n572_), .A3(new_n362_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n361_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n571_), .A2(new_n573_), .A3(KEYINPUT27), .A4(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n493_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n568_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n561_), .A2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n356_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n343_), .A2(new_n262_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n332_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n341_), .B1(new_n583_), .B2(new_n340_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n330_), .A2(new_n331_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n324_), .B1(new_n585_), .B2(KEYINPUT11), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n235_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n581_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT67), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT66), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n343_), .B2(new_n262_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n592_), .A2(new_n593_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n587_), .B2(new_n235_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n343_), .A2(new_n262_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n595_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n591_), .B1(new_n600_), .B2(new_n581_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n599_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n587_), .A2(new_n235_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n603_));
  AND4_X1   g402(.A1(new_n591_), .A2(new_n602_), .A3(new_n581_), .A4(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n590_), .B1(new_n601_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  NAND2_X1  g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n587_), .A2(new_n235_), .A3(new_n596_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n598_), .B1(new_n343_), .B2(new_n262_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n581_), .B(new_n603_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT67), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n602_), .A2(new_n591_), .A3(new_n581_), .A4(new_n603_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n610_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n590_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n611_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(KEYINPUT13), .A3(new_n619_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n321_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n252_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n272_), .A2(new_n321_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT81), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n628_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n263_), .A2(new_n266_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n635_), .B2(new_n626_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n633_), .B1(new_n636_), .B2(new_n631_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n632_), .B1(new_n637_), .B2(KEYINPUT81), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G169gat), .B(G197gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n638_), .B(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n625_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n580_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n316_), .A3(new_n493_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT38), .ZN(new_n649_));
  INV_X1    g448(.A(new_n354_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n625_), .A2(new_n644_), .A3(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT99), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n304_), .A2(new_n305_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n561_), .B2(new_n578_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(KEYINPUT99), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n577_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n649_), .A2(new_n657_), .ZN(G1324gat));
  INV_X1    g457(.A(new_n576_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n647_), .A2(new_n317_), .A3(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n656_), .A2(new_n576_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G8gat), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT100), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n663_), .A2(new_n664_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n664_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n660_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT40), .B(new_n660_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n656_), .B2(new_n521_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT41), .Z(new_n675_));
  OR2_X1    g474(.A1(new_n521_), .A2(G15gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n646_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT101), .ZN(G1326gat));
  OAI21_X1  g477(.A(G22gat), .B1(new_n656_), .B2(new_n560_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT42), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n560_), .A2(G22gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n646_), .B2(new_n681_), .ZN(G1327gat));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n568_), .A2(new_n577_), .A3(new_n576_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n520_), .B(new_n559_), .C1(new_n486_), .C2(new_n499_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n292_), .A2(new_n302_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT79), .B1(new_n687_), .B2(KEYINPUT37), .ZN(new_n688_));
  INV_X1    g487(.A(new_n306_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n312_), .B2(new_n202_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n690_), .B2(KEYINPUT79), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n561_), .A2(new_n578_), .A3(KEYINPUT103), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n686_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT43), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n691_), .A2(new_n695_), .A3(new_n579_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT104), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n691_), .A2(new_n698_), .A3(new_n695_), .A4(new_n579_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n694_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n625_), .A2(new_n644_), .A3(new_n354_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT102), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n700_), .B2(new_n702_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n577_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n653_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n561_), .B2(new_n578_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n701_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n493_), .A2(new_n241_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT105), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n706_), .A2(new_n241_), .B1(new_n710_), .B2(new_n712_), .ZN(G1328gat));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n243_), .A3(new_n659_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT45), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n700_), .A2(new_n702_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n720_), .A2(KEYINPUT106), .A3(new_n659_), .A4(new_n703_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(G36gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n659_), .A3(new_n703_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n716_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT46), .B(new_n717_), .C1(new_n722_), .C2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n724_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n728_), .A2(KEYINPUT107), .A3(G36gat), .A4(new_n721_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n717_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n726_), .A2(new_n731_), .ZN(G1329gat));
  NAND4_X1  g531(.A1(new_n720_), .A2(G43gat), .A3(new_n520_), .A4(new_n703_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n710_), .A2(new_n521_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(G43gat), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g535(.A1(new_n709_), .A2(new_n542_), .A3(new_n559_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n704_), .A2(new_n705_), .A3(new_n560_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(new_n542_), .ZN(G1331gat));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n624_), .A2(new_n643_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n580_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n742_), .B2(new_n577_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT108), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n654_), .A2(new_n354_), .A3(new_n741_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n745_), .A2(new_n740_), .A3(new_n577_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1332gat));
  OAI21_X1  g546(.A(G64gat), .B1(new_n745_), .B2(new_n576_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT48), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n576_), .A2(G64gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n742_), .B2(new_n750_), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n745_), .B2(new_n521_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT49), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n520_), .A2(new_n325_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n742_), .B2(new_n754_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n745_), .B2(new_n560_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n559_), .A2(new_n329_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n742_), .B2(new_n758_), .ZN(G1335gat));
  AND3_X1   g558(.A1(new_n708_), .A2(new_n650_), .A3(new_n741_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n493_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n700_), .A2(new_n650_), .A3(new_n741_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n577_), .A2(new_n203_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(G1336gat));
  AOI21_X1  g563(.A(G92gat), .B1(new_n760_), .B2(new_n659_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n576_), .A2(new_n204_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n762_), .B2(new_n766_), .ZN(G1337gat));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n211_), .B1(new_n762_), .B2(new_n520_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n760_), .B(new_n520_), .C1(new_n210_), .C2(new_n212_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n768_), .B1(new_n773_), .B2(KEYINPUT51), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n772_), .A2(KEYINPUT109), .A3(new_n775_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n772_), .A2(KEYINPUT110), .A3(new_n775_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT110), .B1(new_n772_), .B2(new_n775_), .ZN(new_n778_));
  OAI22_X1  g577(.A1(new_n774_), .A2(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n760_), .A2(new_n208_), .A3(new_n559_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n762_), .A2(new_n559_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(G106gat), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT52), .B(new_n208_), .C1(new_n762_), .C2(new_n559_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g585(.A1(new_n314_), .A2(new_n644_), .A3(new_n624_), .A4(new_n354_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT54), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n629_), .A2(new_n630_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n634_), .B(new_n631_), .C1(new_n635_), .C2(new_n626_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n641_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n638_), .B2(new_n642_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n603_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n581_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n602_), .A2(KEYINPUT111), .A3(new_n603_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n601_), .B2(new_n604_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n795_), .A2(KEYINPUT112), .A3(new_n796_), .A4(new_n797_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n600_), .A2(KEYINPUT55), .A3(new_n581_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n610_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n619_), .B(new_n792_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n589_), .B(new_n610_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n805_), .A2(new_n610_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n792_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n691_), .A2(new_n810_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n643_), .A2(new_n619_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n620_), .B2(new_n792_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n618_), .B1(new_n617_), .B2(new_n590_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n792_), .B(new_n823_), .C1(new_n825_), .C2(new_n811_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n820_), .B(new_n653_), .C1(new_n822_), .C2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n819_), .B1(new_n829_), .B2(KEYINPUT115), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n643_), .A2(new_n619_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n620_), .A2(new_n792_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT113), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n826_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n707_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n820_), .B1(new_n837_), .B2(KEYINPUT57), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n818_), .B1(new_n830_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n788_), .B1(new_n841_), .B2(new_n354_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n659_), .A2(new_n577_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n567_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n643_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n841_), .B2(new_n354_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n837_), .B1(new_n836_), .B2(new_n820_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n852_), .A2(new_n819_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT116), .B(new_n650_), .C1(new_n853_), .C2(new_n818_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n788_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n845_), .A2(KEYINPUT59), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n847_), .A2(KEYINPUT59), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n857_), .A2(KEYINPUT117), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT117), .B1(new_n857_), .B2(new_n858_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n643_), .A2(G113gat), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT118), .Z(new_n863_));
  AOI21_X1  g662(.A(new_n849_), .B1(new_n861_), .B2(new_n863_), .ZN(G1340gat));
  NOR2_X1   g663(.A1(new_n624_), .A2(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n848_), .B1(KEYINPUT60), .B2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n866_), .A2(new_n625_), .A3(new_n857_), .A4(new_n858_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(KEYINPUT60), .B2(new_n866_), .ZN(G1341gat));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n848_), .A2(new_n870_), .A3(new_n354_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n859_), .A2(new_n860_), .A3(new_n650_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n870_), .ZN(G1342gat));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n848_), .A2(new_n874_), .A3(new_n653_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n859_), .A2(new_n860_), .A3(new_n314_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n874_), .ZN(G1343gat));
  INV_X1    g676(.A(new_n562_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n842_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n843_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n644_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT119), .B(G141gat), .Z(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1344gat));
  INV_X1    g682(.A(new_n880_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n625_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n880_), .A2(new_n650_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT61), .B(G155gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  AND3_X1   g688(.A1(new_n884_), .A2(G162gat), .A3(new_n691_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G162gat), .B1(new_n884_), .B2(new_n653_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1347gat));
  NOR2_X1   g691(.A1(new_n576_), .A2(new_n493_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n844_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n855_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n643_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G169gat), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT120), .B(KEYINPUT62), .Z(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n896_), .A2(new_n398_), .A3(new_n643_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n897_), .A2(G169gat), .A3(new_n899_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(G1348gat));
  AOI21_X1  g703(.A(G176gat), .B1(new_n896_), .B2(new_n625_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n842_), .A2(new_n895_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n624_), .A2(new_n399_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  AOI21_X1  g707(.A(G183gat), .B1(new_n906_), .B2(new_n354_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n650_), .A2(new_n380_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n896_), .B2(new_n910_), .ZN(G1350gat));
  NAND3_X1  g710(.A1(new_n896_), .A2(new_n653_), .A3(new_n382_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n896_), .A2(new_n691_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(G190gat), .ZN(new_n915_));
  AOI211_X1 g714(.A(KEYINPUT121), .B(new_n386_), .C1(new_n896_), .C2(new_n691_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n912_), .B1(new_n915_), .B2(new_n916_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n879_), .A2(new_n643_), .A3(new_n893_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n918_), .A2(KEYINPUT122), .A3(new_n364_), .ZN(new_n919_));
  AOI21_X1  g718(.A(KEYINPUT122), .B1(new_n918_), .B2(new_n364_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n364_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(G1352gat));
  NAND3_X1  g721(.A1(new_n842_), .A2(new_n878_), .A3(new_n893_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n624_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n367_), .A2(KEYINPUT123), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n924_), .B(new_n925_), .Z(G1353gat));
  NOR2_X1   g725(.A1(new_n923_), .A2(new_n650_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n929_), .A3(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT124), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n927_), .A2(new_n933_), .A3(new_n929_), .A4(new_n930_), .ZN(new_n934_));
  OR3_X1    g733(.A1(new_n927_), .A2(KEYINPUT125), .A3(new_n929_), .ZN(new_n935_));
  OAI21_X1  g734(.A(KEYINPUT125), .B1(new_n927_), .B2(new_n929_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n932_), .A2(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  XNOR2_X1  g736(.A(KEYINPUT127), .B(G218gat), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n923_), .A2(new_n314_), .A3(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n923_), .A2(new_n707_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n940_), .B(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n939_), .B1(new_n942_), .B2(new_n938_), .ZN(G1355gat));
endmodule


