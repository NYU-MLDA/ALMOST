//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT18), .B(G64gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT23), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT80), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT23), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(new_n219_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n212_), .A2(KEYINPUT79), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n212_), .A2(KEYINPUT79), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n215_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT24), .B1(new_n218_), .B2(new_n219_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  MUX2_X1   g027(.A(new_n227_), .B(KEYINPUT24), .S(new_n228_), .Z(new_n229_));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT26), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n231_), .B(new_n232_), .Z(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT25), .B(G183gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(new_n230_), .B2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n226_), .B(new_n229_), .C1(new_n233_), .C2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n223_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT88), .B(G197gat), .ZN(new_n240_));
  MUX2_X1   g039(.A(new_n239_), .B(new_n240_), .S(G204gat), .Z(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G204gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(G197gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT89), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n240_), .A2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT21), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G211gat), .B(G218gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT90), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n250_), .A2(new_n242_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(new_n241_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT20), .B1(new_n238_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n226_), .B1(G183gat), .B2(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n222_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n234_), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT26), .B(G190gat), .Z(new_n258_));
  OAI211_X1 g057(.A(new_n216_), .B(new_n229_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n253_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n254_), .B1(KEYINPUT94), .B2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(KEYINPUT94), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n209_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n238_), .A2(new_n253_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n266_), .B(KEYINPUT20), .C1(new_n253_), .C2(new_n260_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(new_n208_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n206_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(KEYINPUT94), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n270_), .B(KEYINPUT20), .C1(new_n253_), .C2(new_n238_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n208_), .B1(new_n271_), .B2(new_n263_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n268_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n206_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT95), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n269_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n265_), .A2(new_n268_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(KEYINPUT95), .A3(new_n274_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n262_), .A2(new_n209_), .A3(new_n264_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n267_), .A2(new_n208_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n206_), .B(KEYINPUT98), .ZN(new_n285_));
  OAI211_X1 g084(.A(KEYINPUT27), .B(new_n275_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT96), .Z(new_n289_));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT84), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(G155gat), .B2(G162gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n293_), .B(KEYINPUT86), .C1(G155gat), .C2(G162gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT83), .Z(new_n300_));
  OR2_X1    g099(.A1(new_n300_), .A2(KEYINPUT2), .ZN(new_n301_));
  NAND3_X1  g100(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT85), .ZN(new_n303_));
  OR2_X1    g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT3), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(KEYINPUT85), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(KEYINPUT3), .ZN(new_n307_));
  AND4_X1   g106(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n298_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n293_), .B2(KEYINPUT1), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(KEYINPUT1), .B2(new_n293_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n300_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n304_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT82), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n316_), .A2(KEYINPUT97), .A3(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n314_), .A2(new_n304_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n298_), .A2(new_n309_), .B1(new_n313_), .B2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n318_), .B(new_n319_), .Z(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n290_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n323_), .A2(new_n324_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT4), .B1(new_n327_), .B2(KEYINPUT97), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n289_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n325_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(new_n327_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n288_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G1gat), .B(G29gat), .ZN(new_n334_));
  INV_X1    g133(.A(G85gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT0), .B(G57gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  NOR2_X1   g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT30), .B(G43gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT31), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n238_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT81), .B(G15gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n320_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G71gat), .B(G99gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n348_), .B(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n356_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n253_), .B2(KEYINPUT91), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n253_), .B1(new_n323_), .B2(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n367_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT92), .ZN(new_n371_));
  XOR2_X1   g170(.A(G78gat), .B(G106gat), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n371_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n363_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n373_), .A2(KEYINPUT93), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n370_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n370_), .A2(new_n379_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n380_), .B(new_n381_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n353_), .A2(new_n378_), .A3(new_n382_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n287_), .A2(new_n343_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n382_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n281_), .A2(new_n385_), .A3(new_n342_), .A4(new_n286_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n329_), .A2(new_n332_), .A3(KEYINPUT33), .A4(new_n340_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n288_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n340_), .B1(new_n331_), .B2(new_n289_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n277_), .A2(new_n279_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n274_), .A2(KEYINPUT32), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n278_), .B2(new_n396_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n394_), .A2(new_n395_), .B1(new_n343_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n386_), .B1(new_n399_), .B2(new_n385_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n353_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n384_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G71gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT67), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT67), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G71gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n406_), .A3(G78gat), .ZN(new_n407_));
  INV_X1    g206(.A(G57gat), .ZN(new_n408_));
  INV_X1    g207(.A(G64gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT11), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G57gat), .A2(G64gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(G78gat), .B1(new_n404_), .B2(new_n406_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT68), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n415_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT68), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n413_), .A4(new_n407_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n410_), .A2(new_n412_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(new_n411_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n416_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(G106gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(KEYINPUT65), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT7), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT7), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n431_), .A2(new_n427_), .A3(new_n428_), .A4(KEYINPUT65), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n435_), .A2(new_n437_), .A3(KEYINPUT66), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT66), .B1(new_n435_), .B2(new_n437_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n433_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G85gat), .B(G92gat), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT8), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n436_), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n430_), .B(new_n432_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT8), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n441_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n443_), .A2(new_n448_), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n335_), .A2(new_n203_), .A3(KEYINPUT9), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT10), .B(G99gat), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n428_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n441_), .A2(KEYINPUT9), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n451_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT69), .B1(new_n449_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n435_), .A2(new_n437_), .A3(KEYINPUT66), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n430_), .A4(new_n432_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n447_), .B1(new_n460_), .B2(new_n441_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n446_), .A2(new_n447_), .A3(new_n441_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n455_), .B(KEYINPUT69), .C1(new_n461_), .C2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n426_), .B1(new_n456_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n416_), .A2(new_n419_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n421_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n416_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n455_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT12), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n471_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G230gat), .A2(G233gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n475_), .B(KEYINPUT64), .Z(new_n476_));
  NAND3_X1  g275(.A1(new_n465_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n476_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n455_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(new_n424_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n470_), .A2(new_n471_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n478_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G120gat), .B(G148gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(new_n244_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT5), .B(G176gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n477_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT13), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(KEYINPUT13), .A3(new_n491_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT70), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G29gat), .B(G36gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n498_), .B(KEYINPUT70), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n501_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507_));
  INV_X1    g306(.A(G1gat), .ZN(new_n508_));
  INV_X1    g307(.A(G8gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G1gat), .B(G8gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n503_), .A2(new_n505_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT15), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n497_), .B(new_n514_), .C1(new_n516_), .C2(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT75), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n506_), .A2(KEYINPUT15), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT15), .B1(new_n503_), .B2(new_n505_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n513_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT75), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n497_), .A4(new_n514_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n515_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n514_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(G229gat), .A3(G233gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n518_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(G197gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT76), .B(G169gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n518_), .A2(new_n526_), .A3(new_n529_), .A4(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n496_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n402_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n522_), .B1(new_n456_), .B2(new_n464_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT34), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI22_X1  g347(.A1(new_n471_), .A2(new_n515_), .B1(KEYINPUT35), .B2(new_n544_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n542_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n471_), .A2(new_n552_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n553_), .A2(new_n463_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n547_), .B1(new_n554_), .B2(new_n549_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT36), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n551_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n551_), .A2(new_n555_), .A3(KEYINPUT71), .A4(new_n560_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n541_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n558_), .B(KEYINPUT36), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n565_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  AOI221_X4 g370(.A(new_n568_), .B1(new_n541_), .B2(KEYINPUT37), .C1(new_n563_), .C2(new_n564_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n513_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n424_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579_));
  INV_X1    g378(.A(G211gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT16), .B(G183gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  MUX2_X1   g382(.A(new_n576_), .B(new_n578_), .S(new_n583_), .Z(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT17), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n578_), .A2(new_n583_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n586_), .A2(KEYINPUT17), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n573_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT74), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n540_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n342_), .B(KEYINPUT100), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n508_), .A3(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(KEYINPUT101), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(KEYINPUT101), .ZN(new_n597_));
  AND2_X1   g396(.A1(KEYINPUT102), .A2(KEYINPUT38), .ZN(new_n598_));
  NOR2_X1   g397(.A1(KEYINPUT102), .A2(KEYINPUT38), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n596_), .B(new_n597_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n589_), .A2(new_n569_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n540_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n602_), .B2(new_n342_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT103), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n596_), .A2(new_n597_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n600_), .B(new_n604_), .C1(new_n605_), .C2(new_n598_), .ZN(G1324gat));
  NAND3_X1  g405(.A1(new_n540_), .A2(new_n287_), .A3(new_n601_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G8gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT39), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n592_), .A2(new_n509_), .A3(new_n287_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n609_), .A2(KEYINPUT40), .A3(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1325gat));
  OAI21_X1  g414(.A(G15gat), .B1(new_n602_), .B2(new_n401_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT41), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(KEYINPUT41), .ZN(new_n618_));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n592_), .A2(new_n619_), .A3(new_n353_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(G1326gat));
  INV_X1    g422(.A(new_n385_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G22gat), .B1(new_n602_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT42), .ZN(new_n626_));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n592_), .A2(new_n627_), .A3(new_n385_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1327gat));
  INV_X1    g428(.A(new_n573_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT43), .B1(new_n402_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n343_), .A2(new_n398_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n393_), .B1(new_n279_), .B2(new_n277_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n624_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n353_), .B1(new_n635_), .B2(new_n386_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n632_), .B(new_n573_), .C1(new_n636_), .C2(new_n384_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n631_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n589_), .A2(new_n496_), .A3(new_n538_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n639_), .A2(new_n640_), .B1(KEYINPUT107), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n638_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT107), .B1(new_n642_), .B2(KEYINPUT106), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n647_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n638_), .A2(new_n649_), .A3(new_n645_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n593_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(G29gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n569_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n588_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n540_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n343_), .A2(new_n652_), .ZN(new_n656_));
  OAI22_X1  g455(.A1(new_n651_), .A2(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n287_), .A2(KEYINPUT108), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n287_), .A2(KEYINPUT108), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AND4_X1   g460(.A1(new_n658_), .A2(new_n540_), .A3(new_n654_), .A4(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n287_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n666_), .B2(new_n658_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n664_), .B(new_n668_), .C1(new_n666_), .C2(new_n658_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1329gat));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n649_), .B1(new_n638_), .B2(new_n645_), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n647_), .B(new_n644_), .C1(new_n631_), .C2(new_n637_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n353_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G43gat), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n655_), .A2(G43gat), .A3(new_n401_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n673_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT47), .B(new_n678_), .C1(new_n676_), .C2(G43gat), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1330gat));
  INV_X1    g481(.A(G50gat), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n648_), .A2(new_n650_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(new_n385_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n385_), .A2(new_n683_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n655_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT110), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n624_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n690_));
  OAI221_X1 g489(.A(new_n689_), .B1(new_n655_), .B2(new_n686_), .C1(new_n690_), .C2(new_n683_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(G1331gat));
  NOR3_X1   g491(.A1(new_n402_), .A2(new_n538_), .A3(new_n496_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(new_n591_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n594_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n601_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n696_), .A2(new_n408_), .A3(new_n342_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1332gat));
  INV_X1    g497(.A(new_n661_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G64gat), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT48), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n694_), .A2(new_n409_), .A3(new_n661_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1333gat));
  OAI21_X1  g502(.A(G71gat), .B1(new_n696_), .B2(new_n401_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n694_), .A2(new_n403_), .A3(new_n353_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1334gat));
  OAI21_X1  g507(.A(G78gat), .B1(new_n696_), .B2(new_n624_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT50), .ZN(new_n710_));
  INV_X1    g509(.A(G78gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n694_), .A2(new_n711_), .A3(new_n385_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1335gat));
  NAND2_X1  g512(.A1(new_n693_), .A2(new_n654_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n335_), .B1(new_n714_), .B2(new_n593_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n496_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n538_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n589_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n631_), .B2(new_n637_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n343_), .A2(G85gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT112), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n715_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT113), .Z(G1336gat));
  INV_X1    g523(.A(new_n714_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G92gat), .B1(new_n725_), .B2(new_n287_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n699_), .A2(new_n203_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n719_), .B2(new_n727_), .ZN(G1337gat));
  OAI21_X1  g527(.A(G99gat), .B1(new_n720_), .B2(new_n401_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n725_), .A2(new_n452_), .A3(new_n353_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n725_), .A2(new_n428_), .A3(new_n385_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n719_), .A2(new_n385_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G106gat), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT52), .B(new_n428_), .C1(new_n719_), .C2(new_n385_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n734_), .B(new_n740_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(KEYINPUT119), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n465_), .A2(new_n474_), .A3(new_n746_), .A4(new_n476_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n489_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n425_), .B1(new_n480_), .B2(new_n424_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n481_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n470_), .A2(KEYINPUT12), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n553_), .B2(new_n463_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n478_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(KEYINPUT55), .A3(new_n477_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n748_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n748_), .B2(new_n754_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n491_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n534_), .B1(new_n528_), .B2(new_n497_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n514_), .B1(new_n516_), .B2(new_n513_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n761_), .B(new_n762_), .C1(new_n763_), .C2(new_n497_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n497_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT116), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n537_), .A2(new_n764_), .A3(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n759_), .A2(new_n760_), .A3(KEYINPUT58), .A4(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n465_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n476_), .B1(new_n465_), .B2(new_n474_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n746_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n747_), .A2(new_n489_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n748_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(new_n767_), .A3(new_n491_), .A4(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT117), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n776_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n573_), .A2(new_n768_), .A3(new_n777_), .A4(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n773_), .A2(new_n538_), .A3(new_n491_), .A4(new_n774_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n767_), .A2(new_n492_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT57), .B1(new_n782_), .B2(new_n653_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n785_), .B(new_n569_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n779_), .A2(new_n784_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n589_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n717_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n588_), .B(new_n790_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT54), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(KEYINPUT118), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n783_), .A2(new_n786_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n588_), .B1(new_n795_), .B2(new_n779_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n791_), .B(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n593_), .A2(new_n287_), .A3(new_n383_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n793_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n801_), .A2(G113gat), .A3(new_n717_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n789_), .A2(new_n792_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n800_), .A2(new_n805_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n801_), .A2(KEYINPUT59), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n538_), .ZN(new_n808_));
  INV_X1    g607(.A(G113gat), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n745_), .B(new_n803_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n807_), .B2(new_n538_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT119), .B1(new_n811_), .B2(new_n802_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1340gat));
  INV_X1    g612(.A(new_n801_), .ZN(new_n814_));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(KEYINPUT60), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n496_), .B2(KEYINPUT60), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(KEYINPUT120), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n814_), .B(new_n818_), .C1(KEYINPUT120), .C2(new_n817_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n807_), .A2(new_n716_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n815_), .ZN(G1341gat));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n801_), .A2(KEYINPUT59), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n804_), .A2(new_n806_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n588_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G127gat), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n589_), .A2(G127gat), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n801_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n822_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n830_));
  AOI211_X1 g629(.A(KEYINPUT121), .B(new_n828_), .C1(new_n825_), .C2(G127gat), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n814_), .B2(new_n569_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n573_), .A2(G134gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n807_), .B2(new_n834_), .ZN(G1343gat));
  NOR3_X1   g634(.A1(new_n661_), .A2(new_n624_), .A3(new_n593_), .ZN(new_n836_));
  AND4_X1   g635(.A1(new_n401_), .A2(new_n793_), .A3(new_n799_), .A4(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n538_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n716_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  AND3_X1   g640(.A1(new_n793_), .A2(new_n799_), .A3(new_n401_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n836_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT122), .B1(new_n843_), .B2(new_n589_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n837_), .A2(new_n845_), .A3(new_n588_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n844_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1346gat));
  NAND2_X1  g651(.A1(new_n837_), .A2(new_n569_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  INV_X1    g653(.A(G162gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n854_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n843_), .A2(new_n855_), .A3(new_n630_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(G1347gat));
  NAND3_X1  g659(.A1(new_n661_), .A2(new_n353_), .A3(new_n593_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n385_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n804_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G169gat), .B1(new_n865_), .B2(new_n717_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT62), .B(G169gat), .C1(new_n865_), .C2(new_n717_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n865_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(new_n538_), .A3(new_n221_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n868_), .A2(new_n869_), .A3(new_n871_), .ZN(G1348gat));
  AOI21_X1  g671(.A(G176gat), .B1(new_n870_), .B2(new_n716_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n793_), .A2(new_n799_), .A3(new_n624_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n863_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n496_), .A2(new_n219_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n873_), .B1(new_n878_), .B2(new_n879_), .ZN(G1349gat));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n588_), .A3(new_n877_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n589_), .A2(new_n234_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n881_), .A2(new_n210_), .B1(new_n870_), .B2(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n865_), .B2(new_n630_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n653_), .A2(new_n258_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n865_), .B2(new_n885_), .ZN(G1351gat));
  NOR3_X1   g685(.A1(new_n699_), .A2(new_n343_), .A3(new_n624_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n842_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n717_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n239_), .ZN(G1352gat));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n496_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n244_), .ZN(G1353gat));
  AOI21_X1  g691(.A(new_n589_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n842_), .A2(new_n887_), .A3(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT126), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n894_), .B(new_n896_), .ZN(G1354gat));
  INV_X1    g696(.A(G218gat), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n888_), .A2(new_n898_), .A3(new_n630_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n842_), .A2(new_n569_), .A3(new_n887_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n900_), .A2(KEYINPUT127), .ZN(new_n901_));
  AOI21_X1  g700(.A(G218gat), .B1(new_n900_), .B2(KEYINPUT127), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n901_), .B2(new_n902_), .ZN(G1355gat));
endmodule


