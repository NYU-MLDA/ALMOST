//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT87), .ZN(new_n203_));
  OR2_X1    g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT85), .B(KEYINPUT2), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n206_), .B(new_n209_), .C1(new_n210_), .C2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT85), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n214_), .B2(KEYINPUT2), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n204_), .B(new_n205_), .C1(new_n213_), .C2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT86), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT83), .B1(new_n205_), .B2(KEYINPUT1), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(G155gat), .A4(G162gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n205_), .A2(KEYINPUT1), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n219_), .A2(new_n222_), .A3(new_n204_), .A4(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n212_), .A2(new_n207_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(KEYINPUT84), .A3(new_n225_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n214_), .A2(KEYINPUT2), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n214_), .A2(KEYINPUT2), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n211_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n233_), .A2(new_n215_), .A3(new_n206_), .A4(new_n209_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT86), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n204_), .A4(new_n205_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n218_), .A2(new_n230_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n203_), .B1(new_n237_), .B2(KEYINPUT29), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT89), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G197gat), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G204gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT88), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n244_), .B2(G204gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT21), .ZN(new_n249_));
  AND2_X1   g048(.A1(G211gat), .A2(G218gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G211gat), .A2(G218gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n246_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT21), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n243_), .A2(new_n245_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n256_), .A2(new_n254_), .A3(KEYINPUT21), .A4(new_n248_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n253_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n238_), .A2(new_n241_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n241_), .B1(new_n238_), .B2(new_n258_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n202_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n218_), .A2(new_n230_), .A3(new_n262_), .A4(new_n236_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G22gat), .B(G50gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT28), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n263_), .A2(new_n265_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT90), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT90), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n266_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n237_), .A2(KEYINPUT29), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(KEYINPUT87), .A3(new_n258_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n240_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n202_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n238_), .A2(new_n241_), .A3(new_n258_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n261_), .A2(new_n273_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n272_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n261_), .B2(new_n279_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n237_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT95), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n237_), .A2(new_n290_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n218_), .A2(new_n230_), .A3(new_n286_), .A4(new_n236_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(KEYINPUT4), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT95), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n237_), .A2(new_n290_), .A3(new_n297_), .A4(new_n291_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n293_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT0), .B(G57gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(G85gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(G1gat), .B(G29gat), .Z(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(KEYINPUT33), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT33), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n303_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(new_n309_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n293_), .A2(new_n296_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT96), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n300_), .A4(new_n298_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT96), .B1(new_n299_), .B2(new_n301_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n294_), .A2(new_n295_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n310_), .B1(new_n319_), .B2(new_n301_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT23), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(G183gat), .A3(G190gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n330_), .A2(KEYINPUT78), .A3(G183gat), .A4(G190gat), .ZN(new_n334_));
  OR2_X1    g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT22), .ZN(new_n339_));
  INV_X1    g138(.A(G176gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AOI211_X1 g140(.A(G169gat), .B(G176gat), .C1(new_n338_), .C2(KEYINPUT22), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n336_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT25), .B(G183gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n329_), .A2(new_n331_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n349_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(KEYINPUT24), .A3(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n347_), .A2(new_n348_), .A3(new_n351_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n344_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n258_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n345_), .A2(new_n346_), .B1(new_n350_), .B2(new_n349_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n353_), .A2(KEYINPUT24), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT91), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT91), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n353_), .A2(new_n361_), .A3(KEYINPUT24), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n352_), .A3(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n358_), .A2(new_n363_), .A3(new_n334_), .A4(new_n333_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n253_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n348_), .A2(new_n335_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT22), .B(G169gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n340_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n353_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT19), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n357_), .A2(new_n370_), .A3(KEYINPUT20), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n362_), .A2(new_n352_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n361_), .B1(new_n353_), .B2(KEYINPUT24), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n334_), .B(new_n333_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n347_), .A2(new_n351_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n369_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n258_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n365_), .A2(new_n344_), .A3(new_n355_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(KEYINPUT20), .A3(new_n381_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(KEYINPUT92), .A2(new_n374_), .B1(new_n382_), .B2(new_n372_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n382_), .A2(KEYINPUT92), .A3(new_n372_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n327_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n374_), .A2(KEYINPUT92), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n372_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(KEYINPUT92), .A3(new_n372_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n326_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT94), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n385_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n388_), .A2(KEYINPUT94), .A3(new_n326_), .A4(new_n389_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n311_), .A2(new_n314_), .A3(new_n321_), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n326_), .A2(KEYINPUT32), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n388_), .A2(new_n389_), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT97), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n357_), .A2(KEYINPUT20), .ZN(new_n399_));
  INV_X1    g198(.A(new_n370_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n372_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT98), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT98), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n403_), .B(new_n372_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n402_), .B(new_n404_), .C1(new_n372_), .C2(new_n382_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(KEYINPUT32), .A3(new_n326_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n313_), .A2(new_n309_), .ZN(new_n407_));
  AOI211_X1 g206(.A(new_n310_), .B(new_n303_), .C1(new_n299_), .C2(new_n301_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n398_), .B(new_n406_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n395_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n305_), .A2(new_n310_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n313_), .A2(new_n309_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n411_), .B(new_n412_), .C1(new_n280_), .C2(new_n282_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n405_), .A2(new_n327_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n415_), .A2(KEYINPUT27), .A3(new_n390_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT27), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n392_), .A2(new_n417_), .A3(new_n393_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT99), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT99), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n392_), .A2(new_n420_), .A3(new_n417_), .A4(new_n393_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n416_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n283_), .A2(new_n410_), .B1(new_n414_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n288_), .A2(KEYINPUT82), .A3(new_n289_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT82), .B1(new_n288_), .B2(new_n289_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT31), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(KEYINPUT31), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT80), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n344_), .A3(new_n355_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n428_), .A2(KEYINPUT80), .A3(new_n356_), .A4(new_n429_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n433_), .B(KEYINPUT79), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT30), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G15gat), .B(G43gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n435_), .B(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n431_), .A2(new_n432_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT100), .B1(new_n423_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n411_), .A2(new_n412_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(new_n283_), .A3(new_n422_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT100), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n419_), .A2(new_n421_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n416_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(new_n413_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n283_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n395_), .B2(new_n409_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n448_), .B(new_n442_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n444_), .A2(new_n447_), .A3(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G85gat), .B(G92gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT7), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G99gat), .A2(G106gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n465_), .B(new_n466_), .C1(new_n459_), .C2(KEYINPUT7), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n458_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT8), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n470_), .B(new_n458_), .C1(new_n462_), .C2(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n457_), .A2(KEYINPUT9), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT9), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  INV_X1    g274(.A(G92gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT64), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n465_), .A2(new_n466_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  INV_X1    g280(.A(G106gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT64), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n473_), .A2(new_n484_), .A3(new_n477_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n479_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G57gat), .B(G64gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT66), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(KEYINPUT11), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G71gat), .A2(G78gat), .ZN(new_n491_));
  OR2_X1    g290(.A1(G71gat), .A2(G78gat), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n491_), .B(new_n492_), .C1(new_n487_), .C2(KEYINPUT11), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n488_), .B1(new_n487_), .B2(KEYINPUT11), .ZN(new_n494_));
  OR3_X1    g293(.A1(new_n490_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n472_), .A2(new_n486_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT67), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT12), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n479_), .A2(new_n485_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n501_), .A2(new_n483_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n495_), .A2(new_n496_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT67), .B(new_n500_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G230gat), .A2(G233gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n503_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n499_), .A2(new_n504_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n497_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n508_), .A2(new_n506_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G120gat), .B(G148gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G176gat), .B(G204gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n510_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT13), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n518_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522_));
  INV_X1    g321(.A(G1gat), .ZN(new_n523_));
  INV_X1    g322(.A(G8gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G8gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT71), .ZN(new_n529_));
  AND2_X1   g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n503_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT16), .B(G183gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G211gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G127gat), .B(G155gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n533_), .B1(KEYINPUT17), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT72), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n539_), .A3(KEYINPUT17), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT73), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n538_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT37), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT69), .B(G43gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G50gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G29gat), .B(G36gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT15), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n472_), .A2(new_n486_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT35), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT70), .B1(new_n502_), .B2(new_n547_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n550_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n553_), .A2(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G134gat), .ZN(new_n561_));
  INV_X1    g360(.A(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n565_));
  INV_X1    g364(.A(new_n558_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n550_), .A2(new_n566_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n559_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n563_), .B(KEYINPUT36), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n559_), .B2(new_n567_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n543_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n559_), .A2(new_n567_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT37), .B(new_n568_), .C1(new_n574_), .C2(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n521_), .A2(new_n542_), .A3(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT74), .ZN(new_n578_));
  INV_X1    g377(.A(new_n528_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n547_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT75), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n548_), .A2(new_n528_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n547_), .A2(new_n579_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n582_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G169gat), .B(G197gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT76), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(G113gat), .ZN(new_n591_));
  INV_X1    g390(.A(G141gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n584_), .A2(new_n587_), .A3(new_n593_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n577_), .B2(KEYINPUT74), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n456_), .A2(new_n578_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n523_), .A3(new_n445_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT38), .ZN(new_n606_));
  INV_X1    g405(.A(new_n542_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n521_), .A2(new_n598_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT102), .B(new_n568_), .C1(new_n574_), .C2(new_n571_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n456_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT103), .B1(new_n456_), .B2(new_n612_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n607_), .B(new_n608_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n445_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n606_), .A2(new_n619_), .ZN(G1324gat));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621_));
  OAI21_X1  g420(.A(G8gat), .B1(new_n617_), .B2(new_n422_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT39), .B(G8gat), .C1(new_n617_), .C2(new_n422_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n602_), .A2(new_n603_), .A3(new_n524_), .A4(new_n451_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT104), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n621_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n627_), .B(new_n630_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n631_), .A2(KEYINPUT40), .A3(new_n625_), .A4(new_n624_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(G1325gat));
  OAI21_X1  g432(.A(G15gat), .B1(new_n617_), .B2(new_n442_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT41), .Z(new_n635_));
  INV_X1    g434(.A(G15gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n604_), .A2(new_n636_), .A3(new_n443_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1326gat));
  OAI21_X1  g437(.A(G22gat), .B1(new_n617_), .B2(new_n283_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT42), .ZN(new_n640_));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n604_), .A2(new_n641_), .A3(new_n453_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(G1327gat));
  NOR2_X1   g442(.A1(new_n607_), .A2(new_n612_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT106), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n456_), .A3(new_n608_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT107), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n645_), .A2(new_n456_), .A3(new_n648_), .A4(new_n608_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n445_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n521_), .A2(new_n607_), .A3(new_n598_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n456_), .A2(new_n653_), .A3(new_n576_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n456_), .B2(new_n576_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n652_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(new_n657_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n456_), .A2(new_n576_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT43), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n456_), .A2(new_n653_), .A3(new_n576_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(new_n658_), .A3(new_n659_), .A4(new_n652_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n618_), .B1(new_n661_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n651_), .B1(new_n667_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n647_), .A2(new_n669_), .A3(new_n451_), .A4(new_n649_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT45), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n422_), .B1(new_n661_), .B2(new_n666_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n669_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n671_), .B(KEYINPUT46), .C1(new_n672_), .C2(new_n669_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  INV_X1    g476(.A(G43gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n661_), .A2(new_n666_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(new_n443_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n650_), .A2(new_n678_), .A3(new_n443_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT47), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n442_), .B1(new_n661_), .B2(new_n666_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n684_), .B(new_n681_), .C1(new_n685_), .C2(new_n678_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n650_), .B2(new_n453_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n283_), .B1(new_n661_), .B2(new_n666_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G50gat), .ZN(G1331gat));
  INV_X1    g489(.A(new_n521_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n597_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n456_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n576_), .A2(new_n542_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n445_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n613_), .B(new_n614_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n607_), .A3(new_n692_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n618_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n699_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g499(.A(G64gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(new_n701_), .A3(new_n451_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n698_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n451_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(G64gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n704_), .B2(G64gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n702_), .B1(new_n707_), .B2(new_n708_), .ZN(G1333gat));
  INV_X1    g508(.A(G71gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n695_), .A2(new_n710_), .A3(new_n443_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n703_), .A2(new_n443_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT49), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(G71gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n712_), .B2(G71gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n715_), .B2(new_n716_), .ZN(G1334gat));
  OAI21_X1  g516(.A(G78gat), .B1(new_n698_), .B2(new_n283_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT50), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n283_), .A2(G78gat), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT108), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n695_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1335gat));
  NAND2_X1  g522(.A1(new_n693_), .A2(new_n645_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n475_), .B1(new_n724_), .B2(new_n618_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT109), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n691_), .A2(new_n607_), .A3(new_n597_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n665_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n618_), .A2(new_n475_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  OAI21_X1  g529(.A(new_n476_), .B1(new_n724_), .B2(new_n422_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT110), .Z(new_n732_));
  NOR2_X1   g531(.A1(new_n422_), .A2(new_n476_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n728_), .B2(new_n733_), .ZN(G1337gat));
  INV_X1    g533(.A(new_n724_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n735_), .A2(new_n481_), .A3(new_n443_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n728_), .A2(new_n443_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G99gat), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(G1338gat));
  OAI211_X1 g539(.A(new_n453_), .B(new_n727_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n665_), .A2(KEYINPUT112), .A3(new_n453_), .A4(new_n727_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(G106gat), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n743_), .A2(new_n744_), .A3(KEYINPUT52), .A4(G106gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n735_), .A2(new_n482_), .A3(new_n453_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n735_), .A2(KEYINPUT111), .A3(new_n482_), .A4(new_n453_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(new_n748_), .A3(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n747_), .A2(new_n756_), .A3(new_n753_), .A4(new_n748_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  NOR2_X1   g557(.A1(new_n451_), .A2(new_n618_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n443_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n453_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(KEYINPUT117), .B2(KEYINPUT59), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n761_), .A2(KEYINPUT117), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n499_), .A2(new_n506_), .A3(new_n504_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT115), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n499_), .A2(new_n504_), .A3(new_n766_), .A4(new_n506_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n765_), .A2(G230gat), .A3(G233gat), .A4(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n507_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT55), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n507_), .A2(new_n769_), .A3(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n768_), .A2(new_n771_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n516_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT56), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n510_), .A2(new_n516_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n581_), .A2(new_n582_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n585_), .A2(new_n583_), .A3(new_n586_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n594_), .A3(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n596_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n774_), .A2(new_n783_), .A3(new_n516_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n776_), .A2(new_n778_), .A3(new_n782_), .A4(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n777_), .B1(new_n775_), .B2(KEYINPUT56), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n782_), .A4(new_n784_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n787_), .A2(new_n576_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n612_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n776_), .A2(new_n597_), .A3(new_n778_), .A4(new_n784_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n782_), .A2(new_n517_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(KEYINPUT57), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n790_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n792_), .A2(new_n793_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n612_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n796_), .A2(KEYINPUT118), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n800_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n787_), .A2(new_n576_), .A3(new_n789_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n607_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n577_), .A2(new_n810_), .A3(new_n598_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n691_), .A2(new_n694_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT54), .B1(new_n814_), .B2(new_n597_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n577_), .A2(KEYINPUT113), .A3(new_n810_), .A4(new_n598_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n762_), .B(new_n763_), .C1(new_n809_), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n760_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n801_), .A2(new_n802_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n607_), .B1(new_n821_), .B2(new_n796_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n283_), .B(new_n820_), .C1(new_n822_), .C2(new_n818_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT59), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n819_), .A2(new_n824_), .A3(G113gat), .A4(new_n597_), .ZN(new_n825_));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n823_), .B2(new_n598_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1340gat));
  NAND3_X1  g627(.A1(new_n819_), .A2(new_n521_), .A3(new_n824_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT119), .B(G120gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n521_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n831_), .B1(new_n823_), .B2(new_n837_), .ZN(G1341gat));
  NOR2_X1   g637(.A1(new_n823_), .A2(new_n542_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(G127gat), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n819_), .A2(new_n824_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n607_), .A2(G127gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(G1342gat));
  INV_X1    g642(.A(new_n576_), .ZN(new_n844_));
  INV_X1    g643(.A(G134gat), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n819_), .A2(new_n824_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n823_), .B2(new_n612_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(KEYINPUT121), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1343gat));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n442_), .B(new_n759_), .C1(new_n822_), .C2(new_n818_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n283_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n794_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT116), .B1(new_n794_), .B2(KEYINPUT57), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n542_), .B1(new_n859_), .B2(new_n806_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n443_), .B1(new_n860_), .B2(new_n817_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n861_), .A2(KEYINPUT122), .A3(new_n453_), .A4(new_n759_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n597_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G141gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n592_), .A3(new_n597_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n863_), .A2(new_n521_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G148gat), .ZN(new_n869_));
  INV_X1    g668(.A(G148gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n863_), .A2(new_n870_), .A3(new_n521_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1345gat));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT123), .Z(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n863_), .B2(new_n607_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n874_), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n542_), .B(new_n876_), .C1(new_n856_), .C2(new_n862_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1346gat));
  AOI21_X1  g677(.A(G162gat), .B1(new_n863_), .B2(new_n791_), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n562_), .B(new_n844_), .C1(new_n856_), .C2(new_n862_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n446_), .A2(new_n451_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n598_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT124), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n283_), .B(new_n884_), .C1(new_n809_), .C2(new_n818_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G169gat), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(KEYINPUT125), .A3(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n804_), .A2(KEYINPUT118), .A3(new_n805_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n808_), .A2(new_n821_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n542_), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n453_), .B(new_n882_), .C1(new_n891_), .C2(new_n817_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n367_), .A3(new_n597_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n887_), .A2(KEYINPUT125), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n887_), .A2(KEYINPUT125), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n885_), .A2(G169gat), .A3(new_n894_), .A4(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n888_), .A2(new_n893_), .A3(new_n896_), .ZN(G1348gat));
  AOI21_X1  g696(.A(G176gat), .B1(new_n892_), .B2(new_n521_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n453_), .B1(new_n860_), .B2(new_n817_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n882_), .A2(new_n691_), .A3(new_n340_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1349gat));
  AOI21_X1  g700(.A(new_n882_), .B1(new_n891_), .B2(new_n817_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n345_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n902_), .A2(new_n607_), .A3(new_n283_), .A4(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n892_), .A2(KEYINPUT126), .A3(new_n607_), .A4(new_n903_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n899_), .A2(new_n607_), .A3(new_n451_), .A4(new_n446_), .ZN(new_n908_));
  INV_X1    g707(.A(G183gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n906_), .A2(new_n907_), .A3(new_n910_), .ZN(G1350gat));
  INV_X1    g710(.A(new_n892_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G190gat), .B1(new_n912_), .B2(new_n844_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n892_), .A2(new_n791_), .A3(new_n346_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1351gat));
  OAI211_X1 g714(.A(new_n442_), .B(new_n414_), .C1(new_n822_), .C2(new_n818_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n422_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n597_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n521_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g720(.A1(new_n861_), .A2(new_n451_), .A3(new_n414_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AND2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n922_), .A2(new_n542_), .A3(new_n923_), .A4(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n917_), .A2(new_n607_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n923_), .ZN(G1354gat));
  NOR3_X1   g726(.A1(new_n922_), .A2(G218gat), .A3(new_n612_), .ZN(new_n928_));
  INV_X1    g727(.A(G218gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n917_), .B2(new_n576_), .ZN(new_n930_));
  OAI21_X1  g729(.A(KEYINPUT127), .B1(new_n928_), .B2(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G218gat), .B1(new_n922_), .B2(new_n844_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n917_), .A2(new_n929_), .A3(new_n791_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n931_), .A2(new_n935_), .ZN(G1355gat));
endmodule


