//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n962_, new_n963_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT73), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT73), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n203_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n203_), .B2(new_n206_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT80), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT80), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215_));
  INV_X1    g014(.A(G1gat), .ZN(new_n216_));
  INV_X1    g015(.A(G8gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT14), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G1gat), .B(G8gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n214_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n211_), .A2(new_n213_), .A3(new_n221_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n229_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n203_), .A2(new_n206_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n207_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n203_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT15), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n221_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n223_), .A2(new_n226_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n228_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G113gat), .B(G141gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G169gat), .B(G197gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n240_), .B(new_n241_), .Z(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n228_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT34), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT35), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G99gat), .A2(G106gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT6), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(G99gat), .A3(G106gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258_));
  OR2_X1    g057(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n259_));
  INV_X1    g058(.A(G106gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n257_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n259_), .A2(KEYINPUT65), .A3(new_n260_), .A4(new_n261_), .ZN(new_n264_));
  INV_X1    g063(.A(G85gat), .ZN(new_n265_));
  INV_X1    g064(.A(G92gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G85gat), .A2(G92gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT9), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT9), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G92gat), .ZN(new_n272_));
  OR2_X1    g071(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n270_), .A2(new_n275_), .A3(KEYINPUT67), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT66), .B(G85gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n272_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n277_), .B1(new_n280_), .B2(new_n269_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n263_), .B(new_n264_), .C1(new_n276_), .C2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT8), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n256_), .A2(KEYINPUT69), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G99gat), .A2(G106gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI22_X1  g087(.A1(KEYINPUT68), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n253_), .A2(new_n255_), .A3(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n284_), .A2(new_n288_), .A3(new_n289_), .A4(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n267_), .A2(new_n268_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n283_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(new_n289_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n283_), .B(new_n294_), .C1(new_n296_), .C2(new_n257_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n282_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n236_), .A2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n210_), .B(new_n282_), .C1(new_n295_), .C2(new_n298_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT76), .B1(new_n249_), .B2(new_n250_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n251_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n236_), .A2(new_n299_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n251_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(KEYINPUT75), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G190gat), .B(G218gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT74), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G134gat), .B(G162gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT36), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n308_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n304_), .A2(KEYINPUT75), .A3(new_n314_), .A4(new_n307_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n304_), .A2(new_n307_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n312_), .A2(new_n313_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n316_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT37), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G127gat), .B(G155gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT16), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G183gat), .B(G211gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT17), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT78), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G231gat), .A2(G233gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n221_), .B(new_n333_), .Z(new_n334_));
  AND2_X1   g133(.A1(G71gat), .A2(G78gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G71gat), .A2(G78gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G57gat), .B(G64gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n338_), .B2(KEYINPUT11), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n338_), .B2(KEYINPUT11), .ZN(new_n341_));
  INV_X1    g140(.A(G64gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G57gat), .ZN(new_n343_));
  INV_X1    g142(.A(G57gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G64gat), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n343_), .A2(new_n345_), .A3(new_n340_), .A4(KEYINPUT11), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n339_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n343_), .A2(new_n345_), .A3(KEYINPUT11), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT70), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n343_), .A2(new_n345_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT11), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n350_), .A2(new_n353_), .A3(new_n337_), .A4(new_n346_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n334_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n332_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n348_), .A2(new_n354_), .A3(KEYINPUT71), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  AOI211_X1 g161(.A(new_n330_), .B(new_n329_), .C1(new_n334_), .C2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n362_), .B2(new_n334_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n321_), .A2(new_n322_), .A3(KEYINPUT37), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n325_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT13), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G120gat), .B(G148gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT5), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G176gat), .B(G204gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n370_), .B(new_n371_), .Z(new_n372_));
  OAI211_X1 g171(.A(new_n282_), .B(new_n355_), .C1(new_n295_), .C2(new_n298_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n360_), .A2(KEYINPUT12), .A3(new_n361_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n262_), .A2(new_n258_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n256_), .A3(new_n264_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT67), .B1(new_n270_), .B2(new_n275_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n280_), .A2(new_n277_), .A3(new_n269_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n253_), .A2(new_n255_), .A3(new_n290_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n290_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n296_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT8), .B1(new_n382_), .B2(new_n293_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n379_), .B1(new_n383_), .B2(new_n297_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n373_), .B1(new_n374_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT12), .B1(new_n299_), .B2(new_n356_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G230gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT64), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n385_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n299_), .A2(new_n356_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n373_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n372_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n386_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n299_), .A2(KEYINPUT12), .A3(new_n361_), .A4(new_n360_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n390_), .A3(new_n373_), .A4(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n392_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n372_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n393_), .A2(KEYINPUT72), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT72), .B1(new_n393_), .B2(new_n399_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n368_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT72), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n389_), .A2(new_n392_), .A3(new_n372_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n398_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(KEYINPUT13), .A3(new_n400_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n367_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n246_), .B1(new_n411_), .B2(KEYINPUT79), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G127gat), .B(G134gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G113gat), .B(G120gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n414_), .A2(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n413_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n414_), .A2(new_n415_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(new_n416_), .A3(KEYINPUT85), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n422_), .B(KEYINPUT31), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G99gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(G71gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT25), .B(G183gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT26), .B(G190gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT24), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(G169gat), .B2(G176gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(G169gat), .B2(G176gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n432_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT23), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(G183gat), .A3(G190gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G183gat), .ZN(new_n441_));
  INV_X1    g240(.A(G190gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT23), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT81), .B(KEYINPUT23), .C1(new_n441_), .C2(new_n442_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n440_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G169gat), .A2(G176gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT22), .B(G169gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT82), .B(G176gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G183gat), .A2(G190gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n443_), .B2(new_n439_), .ZN(new_n453_));
  OAI22_X1  g252(.A1(new_n437_), .A2(new_n447_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT30), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n455_), .A2(new_n456_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n455_), .B(new_n456_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n460_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n428_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n464_), .A3(new_n428_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n424_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n424_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n465_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G8gat), .B(G36gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT18), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G64gat), .B(G92gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G226gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT19), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G211gat), .B(G218gat), .ZN(new_n479_));
  OR2_X1    g278(.A1(G197gat), .A2(G204gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G197gat), .A2(G204gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(KEYINPUT21), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT21), .B1(new_n480_), .B2(new_n481_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n479_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(new_n483_), .B2(new_n479_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n448_), .A2(new_n488_), .A3(KEYINPUT24), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n448_), .B2(KEYINPUT24), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n435_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n429_), .A2(new_n430_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n487_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n490_), .A2(new_n435_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT92), .B(new_n431_), .C1(new_n494_), .C2(new_n489_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n443_), .A2(new_n439_), .B1(new_n432_), .B2(new_n435_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  OAI221_X1 g296(.A(new_n448_), .B1(new_n450_), .B2(new_n449_), .C1(new_n447_), .C2(new_n452_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n486_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n479_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n480_), .A2(new_n481_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT21), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n500_), .B1(new_n503_), .B2(new_n482_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n483_), .A2(new_n479_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT20), .B1(new_n454_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n478_), .B1(new_n499_), .B2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n497_), .A2(new_n486_), .A3(new_n498_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n478_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n454_), .B2(new_n506_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n476_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(new_n476_), .A3(new_n513_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT27), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n476_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n497_), .A2(new_n498_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n507_), .B1(new_n519_), .B2(new_n506_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n510_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n509_), .A2(new_n512_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n478_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n499_), .A2(new_n478_), .A3(new_n507_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(new_n521_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n518_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n516_), .A2(KEYINPUT27), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n517_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G1gat), .B(G29gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT95), .B(G85gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT0), .B(G57gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT86), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G155gat), .A2(G162gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(KEYINPUT1), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT1), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n540_), .A2(KEYINPUT86), .A3(G155gat), .A4(G162gat), .ZN(new_n541_));
  OR2_X1    g340(.A1(G155gat), .A2(G162gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(KEYINPUT1), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n539_), .A2(new_n541_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G141gat), .B(G148gat), .Z(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT3), .ZN(new_n547_));
  INV_X1    g346(.A(G141gat), .ZN(new_n548_));
  INV_X1    g347(.A(G148gat), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .A4(KEYINPUT87), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n551_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G141gat), .A2(G148gat), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT2), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n550_), .A2(new_n552_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n542_), .A2(new_n538_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n546_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT4), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n419_), .A2(new_n560_), .A3(new_n561_), .A4(new_n421_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT94), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G225gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n419_), .A2(new_n560_), .A3(new_n421_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n544_), .A2(new_n545_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n568_), .A3(KEYINPUT4), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n563_), .A2(new_n565_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n568_), .A3(new_n564_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n536_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n562_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n565_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n571_), .B(new_n536_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n572_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT89), .ZN(new_n579_));
  XOR2_X1   g378(.A(G22gat), .B(G50gat), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT29), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n546_), .A2(new_n559_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT28), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT28), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n567_), .A2(new_n585_), .A3(new_n582_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT88), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n584_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n581_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n583_), .A2(KEYINPUT28), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n585_), .B1(new_n567_), .B2(new_n582_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT88), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n584_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n580_), .A3(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n582_), .B1(new_n546_), .B2(new_n559_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G106gat), .B1(new_n486_), .B2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n506_), .B(new_n260_), .C1(new_n582_), .C2(new_n567_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G228gat), .A2(G233gat), .ZN(new_n601_));
  INV_X1    g400(.A(G78gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n579_), .B1(new_n596_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n590_), .A2(new_n595_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n610_), .A2(new_n607_), .A3(KEYINPUT89), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(KEYINPUT90), .A3(new_n607_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT90), .B1(new_n610_), .B2(new_n607_), .ZN(new_n613_));
  OAI22_X1  g412(.A1(new_n609_), .A2(new_n611_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n531_), .A2(new_n578_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n576_), .A2(KEYINPUT33), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n570_), .A2(new_n617_), .A3(new_n571_), .A4(new_n536_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n620_));
  INV_X1    g419(.A(new_n516_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n514_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n515_), .A2(KEYINPUT93), .A3(new_n516_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n563_), .A2(new_n564_), .A3(new_n569_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n536_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n566_), .A2(new_n568_), .A3(new_n565_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n619_), .A2(new_n622_), .A3(new_n623_), .A4(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n476_), .A2(KEYINPUT32), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n508_), .A2(new_n513_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(new_n629_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n630_), .B(new_n632_), .C1(new_n572_), .C2(new_n577_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n614_), .B1(new_n628_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n615_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  AOI211_X1 g435(.A(KEYINPUT97), .B(new_n614_), .C1(new_n633_), .C2(new_n628_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n472_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT98), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n640_), .B(new_n472_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n578_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n472_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n531_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n614_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n639_), .A2(new_n641_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n412_), .B(new_n648_), .C1(KEYINPUT79), .C2(new_n411_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n649_), .A2(new_n216_), .A3(new_n642_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT38), .ZN(new_n651_));
  INV_X1    g450(.A(new_n409_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n246_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n365_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n321_), .B(KEYINPUT99), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n638_), .A2(KEYINPUT98), .B1(new_n645_), .B2(new_n643_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT100), .B(new_n656_), .C1(new_n657_), .C2(new_n641_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659_));
  INV_X1    g458(.A(new_n656_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n647_), .B2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n655_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT101), .B(new_n655_), .C1(new_n658_), .C2(new_n661_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n578_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n651_), .B1(new_n666_), .B2(new_n216_), .ZN(G1324gat));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n647_), .A2(new_n660_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT100), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n647_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n644_), .A3(new_n655_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n217_), .B1(new_n677_), .B2(KEYINPUT39), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT103), .B(new_n668_), .C1(new_n676_), .C2(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n673_), .A2(new_n674_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n668_), .A2(KEYINPUT103), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n681_), .A2(new_n675_), .A3(new_n678_), .A4(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n649_), .A2(new_n217_), .A3(new_n644_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n680_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n680_), .A2(new_n683_), .A3(KEYINPUT40), .A4(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n472_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n649_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT101), .B1(new_n672_), .B2(new_n655_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n665_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n695_), .B2(G15gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n472_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n690_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n692_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT104), .B(new_n692_), .C1(new_n696_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1326gat));
  INV_X1    g503(.A(G22gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n614_), .A2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT105), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n649_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n614_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(new_n705_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(KEYINPUT42), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(KEYINPUT42), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n708_), .B1(new_n712_), .B2(new_n713_), .ZN(G1327gat));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n325_), .A2(new_n366_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT106), .B(new_n715_), .C1(new_n648_), .C2(new_n717_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n715_), .A2(KEYINPUT106), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n647_), .B1(KEYINPUT107), .B2(new_n715_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n721_), .B(new_n716_), .C1(KEYINPUT107), .C2(new_n647_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n653_), .A2(new_n365_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n720_), .A2(KEYINPUT44), .A3(new_n722_), .A4(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n722_), .A2(new_n719_), .A3(new_n718_), .A4(new_n723_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n724_), .A2(new_n727_), .A3(new_n642_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G29gat), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n654_), .A2(new_n321_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n648_), .A2(new_n653_), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n732_), .A2(G29gat), .A3(new_n578_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT108), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n729_), .A2(new_n736_), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1328gat));
  NOR3_X1   g537(.A1(new_n732_), .A2(G36gat), .A3(new_n531_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT45), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n724_), .A2(new_n727_), .A3(new_n644_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G36gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n742_), .A3(KEYINPUT46), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1329gat));
  NAND4_X1  g546(.A1(new_n724_), .A2(new_n727_), .A3(G43gat), .A4(new_n691_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n732_), .A2(new_n472_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(G43gat), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n731_), .B2(new_n614_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n724_), .A2(new_n727_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n614_), .A2(G50gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(G1331gat));
  NOR2_X1   g554(.A1(new_n652_), .A2(new_n367_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT109), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n648_), .A2(new_n757_), .A3(new_n246_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n344_), .A3(new_n642_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n246_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n409_), .A2(new_n760_), .ZN(new_n761_));
  AOI211_X1 g560(.A(new_n654_), .B(new_n761_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n642_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n764_), .B2(new_n344_), .ZN(G1332gat));
  NAND3_X1  g564(.A1(new_n758_), .A2(new_n342_), .A3(new_n644_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n762_), .A2(new_n644_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G64gat), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1333gat));
  NAND3_X1  g570(.A1(new_n758_), .A2(new_n426_), .A3(new_n691_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n762_), .A2(new_n691_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G71gat), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  NAND3_X1  g576(.A1(new_n758_), .A2(new_n602_), .A3(new_n614_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n762_), .A2(new_n614_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G78gat), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT50), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT50), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(G1335gat));
  NOR3_X1   g582(.A1(new_n648_), .A2(new_n730_), .A3(new_n761_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n642_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n720_), .A2(new_n722_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n761_), .A2(new_n365_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n578_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(G1336gat));
  NAND3_X1  g589(.A1(new_n784_), .A2(new_n266_), .A3(new_n644_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n788_), .A2(new_n644_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n266_), .ZN(G1337gat));
  NAND3_X1  g592(.A1(new_n786_), .A2(new_n691_), .A3(new_n787_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G99gat), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n784_), .A2(new_n259_), .A3(new_n261_), .A4(new_n691_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT51), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(new_n799_), .A3(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1338gat));
  NAND3_X1  g600(.A1(new_n784_), .A2(new_n260_), .A3(new_n614_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n720_), .A2(new_n614_), .A3(new_n722_), .A4(new_n787_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n803_), .A2(new_n804_), .A3(G106gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(G106gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT53), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n802_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n410_), .B2(new_n760_), .ZN(new_n813_));
  NOR4_X1   g612(.A1(new_n367_), .A2(new_n409_), .A3(KEYINPUT54), .A4(new_n246_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n223_), .A2(new_n237_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n223_), .A2(KEYINPUT111), .A3(new_n237_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n227_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n242_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n245_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n407_), .B2(new_n400_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n388_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n396_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n385_), .A2(new_n386_), .A3(new_n829_), .A4(new_n388_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n372_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n834_), .B(new_n398_), .C1(new_n828_), .C2(new_n831_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n833_), .A2(new_n835_), .A3(KEYINPUT110), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n405_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n389_), .B1(KEYINPUT55), .B2(new_n826_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n372_), .B1(new_n838_), .B2(new_n830_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n834_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT110), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n837_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n825_), .B1(new_n836_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n321_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(KEYINPUT57), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n246_), .A2(new_n399_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n833_), .B2(KEYINPUT110), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n372_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n840_), .A2(new_n849_), .A3(new_n841_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n824_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n851_), .B2(new_n321_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n823_), .A2(new_n405_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT58), .B(new_n854_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n716_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n840_), .A2(new_n849_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT58), .B1(new_n857_), .B2(new_n854_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n853_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n854_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n862_), .A2(KEYINPUT112), .A3(new_n716_), .A4(new_n855_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n845_), .A2(new_n852_), .A3(new_n859_), .A4(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n815_), .B1(new_n864_), .B2(new_n654_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n691_), .A2(new_n642_), .A3(new_n645_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G113gat), .B1(new_n869_), .B2(new_n246_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n866_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT114), .B(KEYINPUT59), .C1(new_n865_), .C2(new_n866_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n862_), .A2(new_n716_), .A3(new_n855_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n845_), .A2(new_n852_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n815_), .B1(new_n654_), .B2(new_n877_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n866_), .A2(KEYINPUT59), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n875_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n875_), .A2(KEYINPUT115), .A3(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(G113gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n246_), .B2(KEYINPUT116), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(KEYINPUT116), .B2(new_n888_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n870_), .B1(new_n887_), .B2(new_n890_), .ZN(G1340gat));
  OAI21_X1  g690(.A(G120gat), .B1(new_n882_), .B2(new_n652_), .ZN(new_n892_));
  INV_X1    g691(.A(G120gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(new_n652_), .B2(KEYINPUT60), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n869_), .B(new_n894_), .C1(KEYINPUT60), .C2(new_n893_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n892_), .A2(new_n895_), .ZN(G1341gat));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n897_));
  AOI21_X1  g696(.A(KEYINPUT115), .B1(new_n875_), .B2(new_n881_), .ZN(new_n898_));
  AOI211_X1 g697(.A(new_n883_), .B(new_n880_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n365_), .A2(G127gat), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n898_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G127gat), .B1(new_n869_), .B2(new_n365_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n897_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n902_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT117), .B(new_n904_), .C1(new_n886_), .C2(new_n900_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1342gat));
  OAI21_X1  g705(.A(G134gat), .B1(new_n886_), .B2(new_n717_), .ZN(new_n907_));
  INV_X1    g706(.A(G134gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n869_), .A2(new_n908_), .A3(new_n656_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1343gat));
  INV_X1    g709(.A(new_n865_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n691_), .A2(new_n578_), .A3(new_n709_), .A4(new_n644_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n760_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT118), .B(G141gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1344gat));
  NOR2_X1   g715(.A1(new_n913_), .A2(new_n652_), .ZN(new_n917_));
  XOR2_X1   g716(.A(KEYINPUT119), .B(G148gat), .Z(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1345gat));
  NOR2_X1   g718(.A1(new_n913_), .A2(new_n654_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT61), .B(G155gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1346gat));
  INV_X1    g721(.A(new_n913_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G162gat), .B1(new_n923_), .B2(new_n656_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n716_), .A2(G162gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT120), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n923_), .B2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT121), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n878_), .A2(new_n614_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n643_), .A2(new_n644_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n246_), .ZN(new_n933_));
  OR3_X1    g732(.A1(new_n930_), .A2(new_n449_), .A3(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  INV_X1    g734(.A(G169gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n933_), .B(KEYINPUT122), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n929_), .A2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n938_), .B2(KEYINPUT123), .ZN(new_n939_));
  AOI21_X1  g738(.A(KEYINPUT123), .B1(new_n929_), .B2(new_n937_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n935_), .B1(new_n939_), .B2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n929_), .A2(new_n937_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944_));
  OAI21_X1  g743(.A(G169gat), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n945_), .A2(KEYINPUT62), .A3(new_n940_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n934_), .B1(new_n942_), .B2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(KEYINPUT124), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n949_), .B(new_n934_), .C1(new_n942_), .C2(new_n946_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n950_), .ZN(G1348gat));
  NOR2_X1   g750(.A1(new_n930_), .A2(new_n931_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n450_), .B1(new_n952_), .B2(new_n409_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n865_), .A2(new_n614_), .ZN(new_n954_));
  AND3_X1   g753(.A1(new_n932_), .A2(G176gat), .A3(new_n409_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n953_), .B1(new_n954_), .B2(new_n955_), .ZN(G1349gat));
  NOR4_X1   g755(.A1(new_n930_), .A2(new_n429_), .A3(new_n654_), .A4(new_n931_), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT125), .Z(new_n958_));
  NOR2_X1   g757(.A1(new_n931_), .A2(new_n654_), .ZN(new_n959_));
  AOI21_X1  g758(.A(G183gat), .B1(new_n954_), .B2(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n958_), .A2(new_n960_), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n952_), .A2(new_n656_), .A3(new_n430_), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n930_), .A2(new_n717_), .A3(new_n931_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n962_), .B1(new_n963_), .B2(new_n442_), .ZN(G1351gat));
  NOR4_X1   g763(.A1(new_n691_), .A2(new_n642_), .A3(new_n709_), .A4(new_n531_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n911_), .A2(new_n965_), .ZN(new_n966_));
  XOR2_X1   g765(.A(new_n966_), .B(KEYINPUT126), .Z(new_n967_));
  INV_X1    g766(.A(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n246_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n409_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g771(.A(KEYINPUT63), .B(G211gat), .C1(new_n968_), .C2(new_n365_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(KEYINPUT63), .B(G211gat), .ZN(new_n974_));
  NOR3_X1   g773(.A1(new_n967_), .A2(new_n654_), .A3(new_n974_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n973_), .A2(new_n975_), .ZN(G1354gat));
  XOR2_X1   g775(.A(KEYINPUT127), .B(G218gat), .Z(new_n977_));
  NOR3_X1   g776(.A1(new_n967_), .A2(new_n717_), .A3(new_n977_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n968_), .A2(new_n656_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n979_), .B2(new_n977_), .ZN(G1355gat));
endmodule


