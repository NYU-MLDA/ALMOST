//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n206_), .A2(KEYINPUT93), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n206_), .B2(KEYINPUT93), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT94), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(KEYINPUT94), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n216_), .B1(KEYINPUT1), .B2(new_n214_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT92), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n220_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n221_), .B(new_n222_), .C1(KEYINPUT1), .C2(new_n214_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n203_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n206_), .A3(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n218_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n228_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n217_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n225_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n230_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n234_), .A3(KEYINPUT4), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n236_), .B(new_n230_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n202_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n202_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(new_n229_), .B2(new_n234_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G1gat), .B(G29gat), .ZN(new_n242_));
  INV_X1    g041(.A(G85gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G57gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT103), .B1(new_n241_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT104), .ZN(new_n249_));
  INV_X1    g048(.A(new_n246_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n235_), .A2(new_n237_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n239_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n240_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(KEYINPUT103), .A3(new_n246_), .A4(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n248_), .A2(new_n249_), .A3(new_n251_), .A4(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n251_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT104), .B1(new_n257_), .B2(new_n247_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT77), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT75), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G57gat), .A2(G64gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G57gat), .A2(G64gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n261_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G57gat), .ZN(new_n266_));
  INV_X1    g065(.A(G64gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT75), .A3(new_n262_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(KEYINPUT74), .A2(G71gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(KEYINPUT74), .A2(G71gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(G78gat), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G78gat), .ZN(new_n276_));
  AND2_X1   g075(.A1(KEYINPUT74), .A2(G71gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(KEYINPUT74), .A2(G71gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n265_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n272_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n281_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT76), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n270_), .A2(new_n271_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT66), .B(G106gat), .Z(new_n292_));
  INV_X1    g091(.A(G99gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT10), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT10), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G99gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n292_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G99gat), .A2(G106gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT70), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT6), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n303_), .A2(new_n305_), .A3(new_n301_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n300_), .A2(KEYINPUT67), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G85gat), .A2(G92gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT9), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G85gat), .A2(G92gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(G85gat), .A2(G92gat), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n316_), .A2(new_n310_), .A3(KEYINPUT68), .ZN(new_n317_));
  INV_X1    g116(.A(G92gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT9), .B1(new_n243_), .B2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n315_), .B(KEYINPUT69), .C1(new_n317_), .C2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT67), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n321_), .B(new_n292_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT69), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n316_), .A2(new_n310_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n319_), .B1(new_n324_), .B2(new_n312_), .ZN(new_n325_));
  NOR4_X1   g124(.A1(new_n316_), .A2(new_n310_), .A3(KEYINPUT68), .A4(KEYINPUT9), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n323_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n309_), .A2(new_n320_), .A3(new_n322_), .A4(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT8), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(KEYINPUT73), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n307_), .A2(new_n308_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G99gat), .A2(G106gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(KEYINPUT71), .A2(KEYINPUT7), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n334_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(KEYINPUT72), .A3(new_n335_), .A4(new_n336_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n332_), .A2(new_n333_), .A3(new_n339_), .A4(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n331_), .B1(new_n342_), .B2(new_n324_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n303_), .A2(new_n305_), .A3(new_n301_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n333_), .B1(new_n344_), .B2(new_n306_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n341_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n331_), .B(new_n324_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n328_), .B1(new_n343_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n260_), .B1(new_n291_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n324_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n330_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n327_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n347_), .A2(new_n352_), .B1(new_n353_), .B2(new_n309_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n285_), .A2(new_n290_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(KEYINPUT77), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n291_), .A2(new_n349_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G230gat), .A2(G233gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT64), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n291_), .B2(new_n349_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT12), .B1(new_n358_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT12), .ZN(new_n368_));
  AOI211_X1 g167(.A(KEYINPUT78), .B(new_n368_), .C1(new_n291_), .C2(new_n349_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n365_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G176gat), .B(G204gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(G120gat), .B(G148gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n362_), .A2(new_n370_), .A3(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(KEYINPUT13), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT13), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT80), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G29gat), .B(G36gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G43gat), .B(G50gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G15gat), .B(G22gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G1gat), .A2(G8gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT14), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G8gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n394_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n392_), .B(KEYINPUT15), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n400_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G229gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n394_), .B(new_n400_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n394_), .A2(new_n400_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n401_), .A2(KEYINPUT87), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n407_), .B1(new_n413_), .B2(new_n406_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT88), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n389_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G141gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G169gat), .B(G197gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT88), .B1(new_n420_), .B2(KEYINPUT89), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n416_), .A2(new_n420_), .B1(new_n421_), .B2(new_n414_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n388_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT27), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT19), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT99), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(G197gat), .A2(G204gat), .ZN(new_n429_));
  INV_X1    g228(.A(G197gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT97), .B(G204gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(G211gat), .B(G218gat), .Z(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n430_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT21), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(G197gat), .B2(G204gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n432_), .A2(KEYINPUT21), .ZN(new_n437_));
  OAI221_X1 g236(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(KEYINPUT21), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT102), .ZN(new_n441_));
  INV_X1    g240(.A(G183gat), .ZN(new_n442_));
  INV_X1    g241(.A(G190gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT23), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT23), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G183gat), .A3(G190gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n441_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n449_), .B(KEYINPUT102), .C1(G183gat), .C2(G190gat), .ZN(new_n453_));
  INV_X1    g252(.A(G169gat), .ZN(new_n454_));
  INV_X1    g253(.A(G176gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G169gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n457_), .B2(new_n455_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(new_n453_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n444_), .A2(new_n448_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G169gat), .A2(G176gat), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n456_), .ZN(new_n464_));
  AOI211_X1 g263(.A(new_n461_), .B(new_n464_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT26), .B(G190gat), .Z(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT25), .B(G183gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT100), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n465_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n440_), .B1(new_n459_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n438_), .A2(new_n439_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(KEYINPUT91), .A2(KEYINPUT22), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n454_), .B1(new_n472_), .B2(new_n455_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n473_), .B1(new_n463_), .B2(new_n472_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n461_), .B2(new_n451_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n456_), .A2(new_n463_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(KEYINPUT24), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n479_), .B2(new_n450_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT20), .B1(new_n471_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n428_), .B1(new_n470_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n459_), .A2(new_n440_), .A3(new_n469_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n471_), .B2(new_n480_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n426_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n483_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G8gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(new_n318_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT18), .B(G64gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n482_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n482_), .B2(new_n487_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n424_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n470_), .A2(new_n481_), .A3(new_n428_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n486_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT27), .B(new_n493_), .C1(new_n499_), .C2(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G233gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n503_), .A2(KEYINPUT96), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(KEYINPUT96), .ZN(new_n505_));
  OAI221_X1 g304(.A(G228gat), .B1(new_n504_), .B2(new_n505_), .C1(new_n440_), .C2(KEYINPUT98), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT29), .B1(new_n232_), .B2(new_n233_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n471_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n508_), .B2(new_n471_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n507_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n510_), .A3(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G22gat), .B(G50gat), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n232_), .A2(new_n233_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT29), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n517_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n517_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n522_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n516_), .A2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n513_), .A2(new_n515_), .A3(new_n525_), .A4(new_n528_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT105), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n502_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n496_), .A2(new_n530_), .A3(new_n531_), .A4(new_n500_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT105), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G71gat), .B(G99gat), .ZN(new_n538_));
  INV_X1    g337(.A(G43gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n480_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G227gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n228_), .B(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT30), .B(G15gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT31), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n543_), .B(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n546_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n537_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n532_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT33), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n251_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n494_), .A2(new_n495_), .ZN(new_n555_));
  OAI211_X1 g354(.A(KEYINPUT33), .B(new_n250_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n229_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n246_), .B(new_n557_), .C1(new_n252_), .C2(new_n239_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .A4(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n257_), .A2(new_n247_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n492_), .A2(KEYINPUT32), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n482_), .A2(new_n487_), .A3(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n499_), .B2(new_n561_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n559_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n552_), .A2(new_n502_), .B1(new_n532_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n549_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n551_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n354_), .A2(new_n392_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n349_), .A2(new_n402_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT34), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT35), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(KEYINPUT83), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n571_), .A2(KEYINPUT35), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n569_), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(KEYINPUT83), .A3(new_n572_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(KEYINPUT83), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n568_), .A2(new_n569_), .A3(new_n578_), .A4(new_n575_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT81), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT36), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n577_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT82), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT37), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n586_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(KEYINPUT84), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT84), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n577_), .A2(new_n594_), .A3(new_n579_), .A4(new_n584_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n590_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n592_), .B1(new_n597_), .B2(new_n591_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n400_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n355_), .B(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G127gat), .B(G155gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(G211gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT16), .B(G183gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT17), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n605_), .A2(KEYINPUT17), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n601_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT85), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n598_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n423_), .A2(new_n567_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT106), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n423_), .A2(new_n567_), .A3(KEYINPUT106), .A4(new_n613_), .ZN(new_n617_));
  AOI211_X1 g416(.A(G1gat), .B(new_n259_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT107), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n567_), .B2(new_n597_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n532_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n258_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n257_), .A2(new_n247_), .A3(KEYINPUT104), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n621_), .B(new_n502_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n564_), .A2(new_n532_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n566_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n537_), .A2(new_n550_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n619_), .B(new_n597_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n620_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n259_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n423_), .A2(new_n610_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(KEYINPUT38), .A2(new_n618_), .B1(new_n633_), .B2(G1gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n618_), .A2(KEYINPUT38), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT108), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n618_), .A2(KEYINPUT108), .A3(KEYINPUT38), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(G1324gat));
  OAI211_X1 g438(.A(new_n501_), .B(new_n632_), .C1(new_n620_), .C2(new_n629_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(new_n641_), .A3(G8gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n640_), .B2(G8gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n616_), .A2(new_n617_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n502_), .A2(G8gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT109), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT109), .ZN(new_n647_));
  INV_X1    g446(.A(new_n645_), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n647_), .B(new_n648_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n649_));
  OAI22_X1  g448(.A1(new_n642_), .A2(new_n643_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI221_X1 g451(.A(KEYINPUT40), .B1(new_n646_), .B2(new_n649_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  OR3_X1    g453(.A1(new_n614_), .A2(G15gat), .A3(new_n549_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n566_), .B(new_n632_), .C1(new_n620_), .C2(new_n629_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(G15gat), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G15gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT111), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT111), .B(new_n655_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  OR3_X1    g463(.A1(new_n614_), .A2(G22gat), .A3(new_n532_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n630_), .A2(new_n621_), .A3(new_n632_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(G22gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G22gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(G29gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n598_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n672_), .B2(KEYINPUT112), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n611_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n672_), .B(new_n675_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n423_), .A4(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n611_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n683_), .A2(KEYINPUT44), .A3(new_n423_), .A4(new_n679_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(new_n631_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT113), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n671_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n686_), .B2(new_n685_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n423_), .A2(new_n567_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n611_), .A2(new_n597_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n671_), .A3(new_n631_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(G1328gat));
  NAND3_X1  g492(.A1(new_n682_), .A2(new_n501_), .A3(new_n684_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n502_), .A2(G36gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n689_), .A2(new_n690_), .A3(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(KEYINPUT46), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1329gat));
  NAND3_X1  g502(.A1(new_n682_), .A2(new_n566_), .A3(new_n684_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G43gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n691_), .A2(new_n539_), .A3(new_n566_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n705_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1330gat));
  INV_X1    g511(.A(G50gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n691_), .A2(new_n713_), .A3(new_n621_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n682_), .A2(new_n621_), .A3(new_n684_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT115), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n715_), .B2(G50gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1331gat));
  INV_X1    g518(.A(new_n388_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n422_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(new_n567_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n613_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n631_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n722_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n678_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n630_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n259_), .A2(new_n266_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1332gat));
  NAND3_X1  g529(.A1(new_n724_), .A2(new_n267_), .A3(new_n501_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n630_), .A2(new_n501_), .A3(new_n727_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G64gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G64gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n724_), .A2(new_n737_), .A3(new_n566_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n630_), .A2(new_n566_), .A3(new_n727_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(G71gat), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n739_), .B2(G71gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1334gat));
  NAND3_X1  g542(.A1(new_n724_), .A2(new_n276_), .A3(new_n621_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n630_), .A2(new_n621_), .A3(new_n727_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G78gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G78gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1335gat));
  AND2_X1   g548(.A1(new_n723_), .A2(new_n690_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n631_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n683_), .A2(new_n679_), .A3(new_n722_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n259_), .A2(new_n243_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n752_), .B2(new_n753_), .ZN(G1336gat));
  AOI21_X1  g553(.A(G92gat), .B1(new_n750_), .B2(new_n501_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n502_), .A2(new_n318_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n752_), .B2(new_n756_), .ZN(G1337gat));
  NAND2_X1  g556(.A1(new_n752_), .A2(new_n566_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G99gat), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n750_), .B(new_n566_), .C1(new_n299_), .C2(new_n298_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT51), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n760_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1338gat));
  AND2_X1   g564(.A1(new_n621_), .A2(new_n292_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n722_), .A2(new_n567_), .A3(new_n690_), .A4(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT117), .Z(new_n768_));
  NAND4_X1  g567(.A1(new_n683_), .A2(new_n621_), .A3(new_n679_), .A4(new_n722_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n768_), .B(new_n775_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n366_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n368_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n358_), .A2(new_n366_), .A3(KEYINPUT12), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n780_), .A2(new_n781_), .B1(new_n350_), .B2(new_n356_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n364_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n783_));
  OAI22_X1  g582(.A1(new_n782_), .A2(new_n363_), .B1(new_n783_), .B2(KEYINPUT55), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n370_), .A2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n778_), .B(new_n377_), .C1(new_n784_), .C2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n379_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n357_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n361_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n370_), .A2(new_n785_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n783_), .A2(KEYINPUT55), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n778_), .B1(new_n793_), .B2(new_n377_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n788_), .A2(new_n422_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n410_), .A2(new_n412_), .A3(new_n405_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n404_), .A2(new_n406_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n420_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n420_), .B2(new_n414_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n380_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n597_), .B1(new_n795_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT57), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n377_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT56), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n805_), .A2(new_n721_), .A3(new_n379_), .A4(new_n787_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n800_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n597_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n803_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n805_), .A2(new_n379_), .A3(new_n799_), .A4(new_n787_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n598_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n788_), .A2(new_n794_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n799_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n610_), .B1(new_n810_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n422_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OR3_X1    g621(.A1(new_n612_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n612_), .B2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n819_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n631_), .A2(new_n537_), .A3(new_n566_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n721_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n808_), .B1(new_n807_), .B2(new_n597_), .ZN(new_n831_));
  AOI211_X1 g630(.A(KEYINPUT57), .B(new_n596_), .C1(new_n806_), .C2(new_n800_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n818_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n825_), .B1(new_n833_), .B2(new_n678_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n827_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n830_), .ZN(new_n836_));
  OAI22_X1  g635(.A1(new_n828_), .A2(new_n830_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n721_), .A2(G113gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n829_), .B1(new_n838_), .B2(new_n839_), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n837_), .B2(new_n720_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n826_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n835_), .ZN(new_n843_));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n720_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(KEYINPUT60), .B2(new_n844_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n841_), .B1(new_n843_), .B2(new_n846_), .ZN(G1341gat));
  NOR2_X1   g646(.A1(new_n826_), .A2(new_n678_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G127gat), .B1(new_n848_), .B2(new_n835_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n610_), .A2(G127gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n838_), .B2(new_n850_), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n843_), .B2(new_n597_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT120), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n855_), .B(new_n852_), .C1(new_n843_), .C2(new_n597_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n598_), .A2(new_n852_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT121), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n854_), .A2(new_n856_), .B1(new_n838_), .B2(new_n858_), .ZN(G1343gat));
  NAND4_X1  g658(.A1(new_n631_), .A2(new_n621_), .A3(new_n502_), .A4(new_n549_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT122), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n826_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n721_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n388_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n611_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  AOI21_X1  g668(.A(G162gat), .B1(new_n862_), .B2(new_n596_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n672_), .A2(G162gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n862_), .B2(new_n871_), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n621_), .A2(new_n502_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n550_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n834_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n454_), .B1(new_n875_), .B2(new_n721_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT124), .B1(new_n834_), .B2(new_n874_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880_));
  INV_X1    g679(.A(new_n874_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n611_), .B1(new_n810_), .B2(new_n818_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n880_), .B(new_n881_), .C1(new_n882_), .C2(new_n825_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n721_), .A2(new_n457_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT125), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n878_), .B1(new_n884_), .B2(new_n886_), .ZN(G1348gat));
  NAND3_X1  g686(.A1(new_n879_), .A2(new_n883_), .A3(new_n388_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n455_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n842_), .A2(G176gat), .A3(new_n388_), .A4(new_n881_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT126), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n889_), .A2(new_n893_), .A3(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1349gat));
  AOI21_X1  g694(.A(G183gat), .B1(new_n848_), .B2(new_n881_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n884_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n610_), .A2(new_n468_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n884_), .B2(new_n598_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n597_), .A2(new_n466_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n884_), .B2(new_n901_), .ZN(G1351gat));
  NAND3_X1  g701(.A1(new_n552_), .A2(new_n501_), .A3(new_n549_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n826_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n721_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n388_), .ZN(new_n907_));
  MUX2_X1   g706(.A(new_n431_), .B(G204gat), .S(new_n907_), .Z(G1353gat));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n610_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  AND2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n909_), .B2(new_n910_), .ZN(G1354gat));
  AOI21_X1  g712(.A(G218gat), .B1(new_n904_), .B2(new_n596_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n672_), .A2(G218gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n904_), .B2(new_n915_), .ZN(G1355gat));
endmodule


