//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT9), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(G92gat), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT6), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n204_), .A2(new_n207_), .A3(new_n211_), .A4(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n216_), .A2(new_n220_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT68), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n225_));
  OAI22_X1  g024(.A1(new_n224_), .A2(new_n225_), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n216_), .A2(new_n220_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(new_n213_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n202_), .B(KEYINPUT67), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n215_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n213_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n231_), .A2(new_n215_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n214_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G29gat), .B(G36gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(G43gat), .B(G50gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G43gat), .B(G50gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(G29gat), .B(G36gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT15), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G232gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  OAI221_X1 g046(.A(new_n244_), .B1(KEYINPUT35), .B2(new_n247_), .C1(new_n235_), .C2(new_n242_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(KEYINPUT35), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  XNOR2_X1  g049(.A(G190gat), .B(G218gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G134gat), .B(G162gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT36), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n248_), .B(new_n249_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT36), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n253_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT37), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G15gat), .B(G22gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT71), .B(G8gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT14), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G1gat), .ZN(new_n266_));
  INV_X1    g065(.A(G1gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(new_n264_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G8gat), .ZN(new_n270_));
  INV_X1    g069(.A(G8gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(new_n271_), .A3(new_n268_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G231gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G57gat), .B(G64gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT11), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G71gat), .B(G78gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n278_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n277_), .A2(KEYINPUT11), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n280_), .B1(new_n283_), .B2(new_n279_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n276_), .B(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT72), .B(KEYINPUT16), .Z(new_n286_));
  XNOR2_X1  g085(.A(G127gat), .B(G155gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G183gat), .B(G211gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT17), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT17), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n292_), .B1(new_n295_), .B2(new_n285_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n261_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT73), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n235_), .A2(new_n284_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n284_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n300_), .B(new_n214_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(KEYINPUT12), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT12), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n235_), .A2(new_n303_), .A3(new_n284_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G230gat), .A2(G233gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT64), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(new_n301_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT5), .B(G176gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G204gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n316_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n309_), .A2(new_n311_), .A3(new_n318_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n317_), .A2(KEYINPUT13), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT13), .B1(new_n317_), .B2(new_n319_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT69), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n298_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT74), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G229gat), .A2(G233gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n242_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n238_), .A2(new_n241_), .A3(KEYINPUT75), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n273_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n330_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n332_), .A2(KEYINPUT76), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT76), .B1(new_n332_), .B2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n327_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n243_), .A2(new_n273_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n334_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT77), .B1(new_n339_), .B2(new_n327_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n338_), .A2(new_n341_), .A3(new_n326_), .A4(new_n334_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G113gat), .B(G141gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT78), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G169gat), .B(G197gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  NAND4_X1  g145(.A1(new_n337_), .A2(new_n340_), .A3(new_n342_), .A4(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n337_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n346_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n349_), .B(new_n352_), .Z(new_n353_));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT81), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT24), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n355_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n360_), .A2(KEYINPUT80), .A3(G190gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT25), .B(G183gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(G190gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT80), .B1(new_n360_), .B2(G190gat), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n355_), .A2(new_n356_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(G183gat), .A3(G190gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT82), .ZN(new_n369_));
  INV_X1    g168(.A(G183gat), .ZN(new_n370_));
  INV_X1    g169(.A(G190gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT23), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n359_), .A2(new_n365_), .A3(new_n366_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n368_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(G183gat), .B2(G190gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT83), .B(G176gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G169gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n357_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G197gat), .B(G204gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT21), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(KEYINPUT21), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n385_), .A2(new_n382_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT20), .B1(new_n381_), .B2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT90), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n373_), .B1(G183gat), .B2(G190gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n357_), .B(KEYINPUT92), .Z(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n379_), .A3(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n394_));
  OR3_X1    g193(.A1(new_n355_), .A2(new_n358_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT26), .B(G190gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n362_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n354_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n395_), .A2(new_n375_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n388_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT93), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G226gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n390_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n388_), .B(KEYINPUT88), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(new_n393_), .A3(new_n399_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n381_), .B2(new_n388_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n407_), .B1(new_n406_), .B2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n414_));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(KEYINPUT32), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n406_), .B1(new_n390_), .B2(new_n402_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n400_), .A2(new_n388_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n411_), .A3(new_n406_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G57gat), .B(G85gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G155gat), .ZN(new_n431_));
  INV_X1    g230(.A(G162gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n431_), .A2(new_n432_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT1), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n436_), .A2(KEYINPUT87), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n435_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(KEYINPUT87), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G141gat), .A2(G148gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n434_), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n443_), .B(KEYINPUT3), .Z(new_n447_));
  XOR2_X1   g246(.A(new_n441_), .B(KEYINPUT2), .Z(new_n448_));
  OAI211_X1 g247(.A(new_n446_), .B(new_n433_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G113gat), .B(G120gat), .ZN(new_n451_));
  INV_X1    g250(.A(G134gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(G127gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT4), .B1(new_n450_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n455_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n455_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n450_), .A2(KEYINPUT95), .A3(new_n455_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n456_), .B1(new_n463_), .B2(KEYINPUT4), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n430_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n468_), .B(new_n430_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n419_), .B(new_n425_), .C1(new_n469_), .C2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT97), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT97), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n470_), .A2(new_n476_), .A3(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n466_), .A2(KEYINPUT33), .A3(new_n430_), .A4(new_n468_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n421_), .A2(new_n418_), .A3(new_n423_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n418_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n423_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n481_), .B1(new_n420_), .B2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n463_), .A2(new_n465_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n430_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n484_), .B(new_n485_), .C1(new_n464_), .C2(new_n467_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n479_), .A2(new_n480_), .A3(new_n483_), .A4(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n472_), .B1(new_n478_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489_));
  INV_X1    g288(.A(G43gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT30), .B(G15gat), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n374_), .A2(new_n380_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n374_), .B2(new_n380_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G227gat), .A2(G233gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n496_), .B(KEYINPUT84), .Z(new_n497_));
  OR3_X1    g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n492_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n455_), .B(KEYINPUT31), .Z(new_n502_));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n503_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n498_), .A2(new_n492_), .A3(new_n499_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n501_), .A2(new_n505_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n505_), .B1(new_n501_), .B2(new_n507_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n450_), .A2(KEYINPUT29), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G228gat), .A2(G233gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n388_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n408_), .B1(KEYINPUT29), .B2(new_n450_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n514_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n515_), .B(new_n520_), .C1(new_n516_), .C2(new_n514_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G22gat), .B(G50gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n450_), .A2(KEYINPUT29), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n524_), .A2(new_n525_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n523_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n523_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n522_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n519_), .A2(new_n532_), .A3(new_n529_), .A4(new_n521_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n488_), .A2(new_n512_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n511_), .A2(new_n536_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n535_), .B(new_n534_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n469_), .A2(new_n471_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n480_), .A2(new_n483_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT27), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n413_), .A2(new_n481_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n480_), .A3(KEYINPUT27), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n540_), .A2(new_n541_), .A3(new_n544_), .A4(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n353_), .B1(new_n537_), .B2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n325_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n541_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n267_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT38), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n322_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n259_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(new_n296_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(G1gat), .B1(new_n560_), .B2(new_n541_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n549_), .A2(KEYINPUT38), .A3(new_n267_), .A4(new_n552_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n561_), .A3(new_n562_), .ZN(G1324gat));
  NAND2_X1  g362(.A1(new_n544_), .A2(new_n546_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(G8gat), .B1(new_n560_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT99), .B(G8gat), .C1(new_n560_), .C2(new_n565_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(KEYINPUT39), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n263_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n325_), .A2(new_n571_), .A3(new_n564_), .A4(new_n548_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT39), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n567_), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n570_), .A2(new_n572_), .A3(KEYINPUT40), .A4(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(G1325gat));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n580_));
  INV_X1    g379(.A(G15gat), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n549_), .A2(new_n580_), .A3(new_n581_), .A4(new_n511_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n325_), .A2(new_n511_), .A3(new_n548_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT100), .B1(new_n583_), .B2(G15gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G15gat), .B1(new_n560_), .B2(new_n512_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT41), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(G1326gat));
  INV_X1    g387(.A(G22gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n536_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n549_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G22gat), .B1(new_n560_), .B2(new_n536_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT42), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(G1327gat));
  NAND2_X1  g393(.A1(new_n558_), .A2(new_n296_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT102), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n557_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n541_), .ZN(new_n598_));
  AOI21_X1  g397(.A(G29gat), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n349_), .B(new_n352_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n322_), .A2(new_n296_), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT101), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT43), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n537_), .A2(new_n547_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n261_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n259_), .B(KEYINPUT37), .ZN(new_n606_));
  AOI211_X1 g405(.A(KEYINPUT43), .B(new_n606_), .C1(new_n537_), .C2(new_n547_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n602_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT44), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(G29gat), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n599_), .B1(new_n613_), .B2(new_n552_), .ZN(G1328gat));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n564_), .A3(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G36gat), .ZN(new_n616_));
  INV_X1    g415(.A(G36gat), .ZN(new_n617_));
  AND4_X1   g416(.A1(new_n617_), .A2(new_n557_), .A3(new_n564_), .A4(new_n596_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT45), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n616_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n616_), .B2(new_n620_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1329gat));
  NAND4_X1  g423(.A1(new_n610_), .A2(G43gat), .A3(new_n511_), .A4(new_n611_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n548_), .A2(new_n511_), .A3(new_n322_), .A4(new_n596_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n490_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT104), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g429(.A(G50gat), .B1(new_n597_), .B2(new_n590_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n590_), .A2(G50gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n612_), .B2(new_n632_), .ZN(G1331gat));
  INV_X1    g432(.A(new_n322_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n600_), .B1(new_n537_), .B2(new_n547_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n298_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(G57gat), .B1(new_n637_), .B2(new_n552_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n323_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n559_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(new_n541_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n638_), .B1(G57gat), .B2(new_n642_), .ZN(G1332gat));
  OR3_X1    g442(.A1(new_n636_), .A2(G64gat), .A3(new_n565_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G64gat), .B1(new_n641_), .B2(new_n565_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT48), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(KEYINPUT48), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n644_), .B1(new_n646_), .B2(new_n647_), .ZN(G1333gat));
  NAND3_X1  g447(.A1(new_n640_), .A2(new_n559_), .A3(new_n511_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(G71gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT49), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n650_), .B1(new_n649_), .B2(G71gat), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n636_), .A2(G71gat), .A3(new_n512_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(G1334gat));
  NAND3_X1  g457(.A1(new_n640_), .A2(new_n559_), .A3(new_n590_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(G78gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT50), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n660_), .B1(new_n659_), .B2(G78gat), .ZN(new_n664_));
  OR3_X1    g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n636_), .A2(G78gat), .A3(new_n536_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(G1335gat));
  AND2_X1   g467(.A1(new_n640_), .A2(new_n596_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G85gat), .B1(new_n669_), .B2(new_n552_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n296_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n600_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n634_), .B(new_n672_), .C1(new_n605_), .C2(new_n607_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT107), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(KEYINPUT107), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n210_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n541_), .B1(new_n677_), .B2(new_n208_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n670_), .B1(new_n676_), .B2(new_n678_), .ZN(G1336gat));
  AOI21_X1  g478(.A(G92gat), .B1(new_n669_), .B2(new_n564_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n564_), .A2(G92gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n676_), .B2(new_n681_), .ZN(G1337gat));
  AND2_X1   g481(.A1(new_n511_), .A2(new_n205_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n669_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n674_), .A2(new_n511_), .A3(new_n675_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G99gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n687_), .B(new_n689_), .ZN(G1338gat));
  OAI21_X1  g489(.A(G106gat), .B1(new_n673_), .B2(new_n536_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT109), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n693_), .B(G106gat), .C1(new_n673_), .C2(new_n536_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(KEYINPUT52), .A3(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n669_), .A2(new_n206_), .A3(new_n590_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT52), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n691_), .A2(KEYINPUT109), .A3(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n696_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT53), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT53), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n695_), .A2(new_n701_), .A3(new_n696_), .A4(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1339gat));
  INV_X1    g502(.A(KEYINPUT55), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n309_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n302_), .A2(new_n307_), .A3(new_n304_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n302_), .A2(KEYINPUT112), .A3(new_n307_), .A4(new_n304_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n305_), .A2(KEYINPUT55), .A3(new_n308_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n705_), .A2(new_n708_), .A3(new_n709_), .A4(new_n710_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n711_), .A2(KEYINPUT56), .A3(new_n316_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT56), .B1(new_n711_), .B2(new_n316_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n600_), .B(new_n319_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT113), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT56), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n708_), .A2(new_n709_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT55), .B1(new_n305_), .B2(new_n308_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n704_), .B(new_n307_), .C1(new_n302_), .C2(new_n304_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n721_), .B2(new_n318_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n711_), .A2(KEYINPUT56), .A3(new_n316_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n724_), .A2(KEYINPUT113), .A3(new_n600_), .A4(new_n319_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n335_), .A2(new_n336_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n346_), .B1(new_n726_), .B2(new_n326_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n326_), .B2(new_n339_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n347_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n317_), .A2(new_n319_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n716_), .A2(new_n725_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n259_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT57), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n724_), .A2(new_n319_), .A3(new_n729_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT58), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n724_), .A2(KEYINPUT58), .A3(new_n319_), .A4(new_n729_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n739_), .A3(new_n261_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT114), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n732_), .A2(KEYINPUT57), .A3(new_n259_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n738_), .A2(new_n739_), .A3(new_n743_), .A4(new_n261_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n735_), .A2(new_n741_), .A3(new_n742_), .A4(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n296_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n353_), .A2(KEYINPUT110), .A3(new_n671_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n600_), .B2(new_n296_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n749_), .A3(new_n322_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n606_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT54), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n606_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n746_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n538_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n551_), .A2(new_n564_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT59), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n742_), .A2(new_n740_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT57), .B1(new_n732_), .B2(new_n259_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n296_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT115), .B(new_n296_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n757_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT59), .ZN(new_n770_));
  INV_X1    g569(.A(new_n760_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n538_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n762_), .A2(G113gat), .A3(new_n600_), .A4(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(G113gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n761_), .B2(new_n353_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1340gat));
  AOI22_X1  g576(.A1(new_n745_), .A2(new_n296_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n778_), .A2(new_n538_), .A3(new_n771_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n773_), .B(new_n639_), .C1(new_n770_), .C2(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT116), .B(G120gat), .Z(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n781_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n322_), .B2(KEYINPUT60), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n779_), .B(new_n784_), .C1(KEYINPUT60), .C2(new_n783_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n785_), .ZN(G1341gat));
  NAND4_X1  g585(.A1(new_n762_), .A2(G127gat), .A3(new_n671_), .A4(new_n773_), .ZN(new_n787_));
  INV_X1    g586(.A(G127gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n761_), .B2(new_n296_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1342gat));
  NOR2_X1   g589(.A1(new_n606_), .A2(new_n452_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n762_), .A2(new_n773_), .A3(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT117), .B(new_n452_), .C1(new_n761_), .C2(new_n259_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  NOR4_X1   g593(.A1(new_n778_), .A2(new_n259_), .A3(new_n538_), .A4(new_n771_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(G134gat), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n792_), .A2(new_n793_), .A3(new_n796_), .ZN(G1343gat));
  NAND3_X1  g596(.A1(new_n760_), .A2(new_n512_), .A3(new_n590_), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT118), .Z(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n746_), .B2(new_n757_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n600_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT119), .B(G141gat), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(G1344gat));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n639_), .ZN(new_n804_));
  XOR2_X1   g603(.A(KEYINPUT120), .B(G148gat), .Z(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(G1345gat));
  XNOR2_X1  g605(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n807_));
  INV_X1    g606(.A(new_n799_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n758_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(G155gat), .B1(new_n809_), .B2(new_n296_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n800_), .A2(new_n431_), .A3(new_n671_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n431_), .B1(new_n800_), .B2(new_n671_), .ZN(new_n813_));
  NOR4_X1   g612(.A1(new_n778_), .A2(new_n799_), .A3(G155gat), .A4(new_n296_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n807_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n812_), .A2(new_n816_), .ZN(G1346gat));
  NOR3_X1   g616(.A1(new_n809_), .A2(new_n432_), .A3(new_n606_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G162gat), .B1(new_n800_), .B2(new_n558_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1347gat));
  AND2_X1   g619(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n769_), .A2(new_n536_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n551_), .A2(new_n564_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n512_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n600_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT122), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(G169gat), .B(new_n821_), .C1(new_n822_), .C2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n769_), .A2(new_n536_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(new_n600_), .A3(new_n378_), .A4(new_n824_), .ZN(new_n830_));
  INV_X1    g629(.A(G169gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n829_), .B2(new_n826_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n828_), .B(new_n830_), .C1(new_n832_), .C2(new_n833_), .ZN(G1348gat));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n634_), .A3(new_n824_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n778_), .A2(new_n538_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n823_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(G176gat), .A3(new_n837_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n835_), .A2(new_n377_), .B1(new_n639_), .B2(new_n838_), .ZN(G1349gat));
  NOR3_X1   g638(.A1(new_n822_), .A2(new_n512_), .A3(new_n823_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n296_), .A2(new_n362_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n836_), .A2(new_n671_), .A3(new_n837_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n840_), .A2(new_n841_), .B1(new_n370_), .B2(new_n842_), .ZN(G1350gat));
  NAND3_X1  g642(.A1(new_n829_), .A2(new_n261_), .A3(new_n824_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G190gat), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n829_), .A2(new_n558_), .A3(new_n396_), .A4(new_n824_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1351gat));
  NOR3_X1   g646(.A1(new_n565_), .A2(new_n598_), .A3(new_n539_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n758_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n353_), .ZN(new_n850_));
  INV_X1    g649(.A(G197gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(KEYINPUT124), .A3(new_n851_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT124), .B(G197gat), .Z(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n850_), .B2(new_n853_), .ZN(G1352gat));
  NOR2_X1   g653(.A1(new_n849_), .A2(new_n323_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT125), .B(G204gat), .Z(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n855_), .B2(new_n858_), .ZN(G1353gat));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n849_), .A2(new_n296_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n860_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n848_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n778_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n671_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT126), .A3(new_n862_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n862_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n864_), .A2(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1354gat));
  NAND3_X1  g670(.A1(new_n866_), .A2(G218gat), .A3(new_n261_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G218gat), .B1(new_n866_), .B2(new_n558_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT127), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT127), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n849_), .A2(new_n259_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n876_), .B(new_n872_), .C1(new_n877_), .C2(G218gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(G1355gat));
endmodule


