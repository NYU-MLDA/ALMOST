//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_;
  INV_X1    g000(.A(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT25), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT25), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G183gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT78), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n210_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n221_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n220_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT79), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n220_), .B(new_n227_), .C1(new_n222_), .C2(new_n224_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n217_), .A2(new_n219_), .A3(new_n226_), .A4(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT81), .B(G176gat), .Z(new_n230_));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT22), .B1(new_n231_), .B2(new_n211_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n230_), .B(new_n232_), .C1(new_n231_), .C2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n237_), .A3(new_n214_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n229_), .A2(KEYINPUT82), .A3(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G99gat), .ZN(new_n244_));
  INV_X1    g043(.A(G43gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G127gat), .B(G134gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(G113gat), .B(G120gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(G15gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT30), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT31), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n251_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n257_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT84), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT1), .ZN(new_n263_));
  OR2_X1    g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n262_), .B1(new_n261_), .B2(KEYINPUT1), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n260_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n268_), .A2(KEYINPUT85), .A3(new_n264_), .A4(new_n263_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n261_), .A2(KEYINPUT1), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AND3_X1   g070(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT86), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT2), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT2), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n279_), .B(new_n280_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n275_), .B(KEYINPUT3), .ZN(new_n282_));
  NAND3_X1  g081(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT87), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n284_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n281_), .A2(new_n282_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n264_), .A2(new_n261_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n250_), .B1(new_n277_), .B2(new_n289_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n271_), .A2(new_n276_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n250_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(KEYINPUT4), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT93), .Z(new_n296_));
  NOR2_X1   g095(.A1(new_n291_), .A2(new_n292_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT94), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT94), .ZN(new_n300_));
  NOR4_X1   g099(.A1(new_n291_), .A2(new_n300_), .A3(KEYINPUT4), .A4(new_n292_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n294_), .B(new_n296_), .C1(new_n299_), .C2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n290_), .A2(new_n293_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n296_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G1gat), .B(G29gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT95), .B(G85gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT0), .B(G57gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n302_), .A2(new_n305_), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n258_), .A2(new_n259_), .A3(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n315_));
  XNOR2_X1  g114(.A(G8gat), .B(G36gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT18), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n322_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  OR3_X1    g125(.A1(new_n321_), .A2(new_n325_), .A3(new_n322_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n225_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n207_), .A2(new_n209_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n203_), .A2(new_n205_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n215_), .B(new_n330_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G169gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n230_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n237_), .A2(new_n214_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n329_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n329_), .A2(new_n335_), .A3(KEYINPUT92), .A4(new_n338_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n341_), .A2(KEYINPUT20), .A3(new_n345_), .A4(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n329_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT89), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n229_), .A2(KEYINPUT82), .A3(new_n238_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT82), .B1(new_n229_), .B2(new_n238_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n328_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n350_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n241_), .A2(new_n329_), .A3(new_n242_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n335_), .A2(new_n338_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n328_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT91), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(KEYINPUT91), .A3(new_n328_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n355_), .A2(new_n357_), .A3(new_n363_), .ZN(new_n364_));
  AOI211_X1 g163(.A(new_n320_), .B(new_n349_), .C1(new_n364_), .C2(new_n344_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n357_), .A2(new_n363_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT89), .B1(new_n356_), .B2(KEYINPUT20), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n344_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n349_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n319_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n315_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n291_), .A2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n373_), .B(KEYINPUT28), .Z(new_n374_));
  OAI21_X1  g173(.A(new_n328_), .B1(new_n291_), .B2(new_n372_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n375_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(G78gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G106gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G22gat), .B(G50gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n376_), .A2(new_n377_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n368_), .A2(new_n319_), .A3(new_n369_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n355_), .A2(new_n345_), .A3(new_n357_), .A4(new_n363_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n339_), .A2(KEYINPUT20), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n344_), .B1(new_n348_), .B2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n388_), .B(KEYINPUT27), .C1(new_n392_), .C2(new_n319_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n371_), .A2(new_n387_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT98), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n371_), .A2(KEYINPUT98), .A3(new_n393_), .A4(new_n387_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n314_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n258_), .A2(new_n259_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n300_), .B1(new_n290_), .B2(KEYINPUT4), .ZN(new_n400_));
  INV_X1    g199(.A(new_n301_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT96), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n294_), .A4(new_n304_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n294_), .B(new_n304_), .C1(new_n299_), .C2(new_n301_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT96), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n310_), .B1(new_n303_), .B2(new_n296_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n302_), .A2(new_n305_), .A3(new_n310_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n302_), .A2(KEYINPUT33), .A3(new_n305_), .A4(new_n310_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n413_), .A2(new_n365_), .A3(new_n370_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n368_), .A2(new_n369_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n416_), .A2(new_n313_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n387_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n387_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(new_n371_), .A3(new_n393_), .A4(new_n313_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n399_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n398_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G141gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G169gat), .B(G197gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G229gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT76), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G29gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G43gat), .B(G50gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT15), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G15gat), .B(G22gat), .ZN(new_n435_));
  INV_X1    g234(.A(G1gat), .ZN(new_n436_));
  INV_X1    g235(.A(G8gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT14), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G8gat), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n440_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n430_), .B1(new_n434_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n433_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT74), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n428_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n433_), .B1(new_n442_), .B2(new_n441_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT75), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n446_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n447_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n427_), .B1(new_n452_), .B2(KEYINPUT77), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT77), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n450_), .A2(new_n446_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(new_n428_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n454_), .B(new_n426_), .C1(new_n456_), .C2(new_n447_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n423_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G231gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n443_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT66), .B(G71gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(new_n379_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G57gat), .B(G64gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n465_), .B(KEYINPUT11), .Z(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(new_n464_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n462_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT73), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G127gat), .B(G155gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT16), .ZN(new_n474_));
  XOR2_X1   g273(.A(G183gat), .B(G211gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT17), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n472_), .B(new_n478_), .ZN(new_n479_));
  OR3_X1    g278(.A1(new_n470_), .A2(KEYINPUT17), .A3(new_n477_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G232gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT34), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(G85gat), .A2(G92gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT9), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n491_), .A2(KEYINPUT64), .A3(new_n490_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT64), .B1(new_n491_), .B2(new_n490_), .ZN(new_n493_));
  OAI221_X1 g292(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT6), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT10), .B(G99gat), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n494_), .B(new_n496_), .C1(G106gat), .C2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT65), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT7), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n496_), .A2(new_n500_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n489_), .A2(new_n491_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n499_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  AOI211_X1 g307(.A(KEYINPUT8), .B(new_n506_), .C1(new_n503_), .C2(new_n496_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n433_), .B(new_n498_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n498_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(KEYINPUT67), .B(new_n498_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n434_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n488_), .B1(new_n512_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G190gat), .B(G218gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G134gat), .B(G162gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT36), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n512_), .A2(new_n488_), .A3(new_n517_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n519_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n522_), .B(KEYINPUT36), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n519_), .B2(new_n524_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT37), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n524_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n526_), .B1(new_n530_), .B2(new_n518_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n519_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT37), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n482_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G176gat), .B(G204gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT70), .ZN(new_n538_));
  XOR2_X1   g337(.A(G120gat), .B(G148gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(KEYINPUT68), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT12), .B1(new_n513_), .B2(new_n469_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n513_), .A2(new_n469_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n515_), .A2(KEYINPUT12), .A3(new_n469_), .A4(new_n516_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n513_), .B(new_n469_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n544_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n550_), .A2(new_n553_), .A3(new_n544_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n536_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n460_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n313_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n436_), .A3(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT99), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT38), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n525_), .A2(new_n528_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n423_), .A2(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n563_), .A2(new_n458_), .A3(new_n482_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(G1gat), .B1(new_n576_), .B2(new_n313_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n568_), .A2(KEYINPUT99), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n568_), .A2(KEYINPUT99), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(KEYINPUT38), .A3(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n571_), .A2(new_n577_), .A3(new_n580_), .ZN(G1324gat));
  NAND2_X1  g380(.A1(new_n371_), .A2(new_n393_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n565_), .A2(G8gat), .A3(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G8gat), .B1(new_n576_), .B2(new_n583_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT39), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT39), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n587_), .B(G8gat), .C1(new_n576_), .C2(new_n583_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n584_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n589_), .B(new_n591_), .ZN(G1325gat));
  INV_X1    g391(.A(new_n399_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G15gat), .B1(new_n576_), .B2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT41), .Z(new_n595_));
  NAND3_X1  g394(.A1(new_n566_), .A2(new_n253_), .A3(new_n399_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1326gat));
  NAND3_X1  g396(.A1(new_n574_), .A2(new_n420_), .A3(new_n575_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT42), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(G22gat), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n598_), .B2(G22gat), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n387_), .A2(G22gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT101), .ZN(new_n604_));
  OAI22_X1  g403(.A1(new_n601_), .A2(new_n602_), .B1(new_n565_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT102), .ZN(G1327gat));
  NAND2_X1  g405(.A1(new_n572_), .A2(new_n482_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n563_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n460_), .A2(new_n608_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n609_), .A2(G29gat), .A3(new_n313_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n562_), .A2(new_n459_), .A3(new_n482_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n529_), .A2(new_n534_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n398_), .B2(new_n422_), .ZN(new_n617_));
  XOR2_X1   g416(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT43), .ZN(new_n620_));
  OAI221_X1 g419(.A(new_n616_), .B1(KEYINPUT104), .B2(new_n620_), .C1(new_n398_), .C2(new_n422_), .ZN(new_n621_));
  AOI211_X1 g420(.A(new_n611_), .B(new_n614_), .C1(new_n619_), .C2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT105), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n619_), .A2(new_n621_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n614_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n624_), .B1(new_n627_), .B2(new_n611_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n614_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n629_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n567_), .B(new_n623_), .C1(new_n628_), .C2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n631_), .A2(new_n632_), .A3(G29gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n631_), .B2(G29gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n610_), .B1(new_n633_), .B2(new_n634_), .ZN(G1328gat));
  INV_X1    g434(.A(KEYINPUT46), .ZN(new_n636_));
  INV_X1    g435(.A(G36gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n627_), .A2(new_n624_), .A3(new_n611_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT105), .B1(new_n629_), .B2(KEYINPUT44), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n622_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n637_), .B1(new_n640_), .B2(new_n582_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n582_), .A2(new_n637_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n609_), .A2(KEYINPUT45), .A3(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT45), .B1(new_n609_), .B2(new_n642_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n636_), .B1(new_n641_), .B2(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n583_), .B(new_n622_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT46), .B(new_n645_), .C1(new_n648_), .C2(new_n637_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1329gat));
  INV_X1    g449(.A(new_n609_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G43gat), .B1(new_n651_), .B2(new_n399_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n593_), .A2(new_n245_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n640_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n653_), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n658_), .B(new_n622_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n659_), .B2(new_n652_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n660_), .ZN(G1330gat));
  AOI21_X1  g460(.A(G50gat), .B1(new_n651_), .B2(new_n420_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n420_), .A2(G50gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n640_), .B2(new_n663_), .ZN(G1331gat));
  INV_X1    g463(.A(G57gat), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n423_), .A2(new_n458_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n563_), .A3(new_n535_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n667_), .B2(new_n313_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT108), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n574_), .A2(new_n458_), .A3(new_n563_), .A4(new_n481_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n670_), .A2(new_n665_), .A3(new_n313_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1332gat));
  OAI21_X1  g471(.A(G64gat), .B1(new_n670_), .B2(new_n583_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT48), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n583_), .A2(G64gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n667_), .B2(new_n675_), .ZN(G1333gat));
  OAI21_X1  g475(.A(G71gat), .B1(new_n670_), .B2(new_n593_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT49), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n593_), .A2(G71gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n667_), .B2(new_n679_), .ZN(G1334gat));
  OAI21_X1  g479(.A(G78gat), .B1(new_n670_), .B2(new_n387_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n420_), .A2(new_n379_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n667_), .B2(new_n684_), .ZN(G1335gat));
  NOR2_X1   g484(.A1(new_n562_), .A2(new_n607_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n666_), .A2(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n687_), .A2(G85gat), .A3(new_n313_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n562_), .A2(new_n459_), .A3(new_n481_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n625_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n567_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n688_), .B1(G85gat), .B2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT110), .Z(G1336gat));
  INV_X1    g492(.A(new_n687_), .ZN(new_n694_));
  INV_X1    g493(.A(G92gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n582_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n690_), .A2(new_n582_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n695_), .ZN(G1337gat));
  INV_X1    g497(.A(G99gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n690_), .B2(new_n399_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n687_), .A2(new_n593_), .A3(new_n497_), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n700_), .A2(new_n701_), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n702_));
  NAND2_X1  g501(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT112), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n702_), .B(new_n704_), .ZN(G1338gat));
  NAND3_X1  g504(.A1(new_n694_), .A2(new_n381_), .A3(new_n420_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n625_), .A2(new_n420_), .A3(new_n689_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT52), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G106gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G106gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g511(.A(KEYINPUT55), .B1(new_n549_), .B2(KEYINPUT115), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n542_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT55), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n552_), .A2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n547_), .A2(new_n548_), .A3(new_n713_), .A4(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n455_), .A2(new_n430_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n429_), .B1(new_n434_), .B2(new_n443_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(new_n446_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n427_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n452_), .B2(new_n427_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n550_), .A2(new_n553_), .A3(new_n542_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n715_), .A2(new_n718_), .A3(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n720_), .A2(new_n727_), .A3(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n731_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n720_), .A2(new_n727_), .A3(new_n733_), .A4(new_n729_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n616_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n719_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT56), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n459_), .A2(KEYINPUT114), .A3(new_n726_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n719_), .A2(new_n736_), .A3(KEYINPUT56), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n726_), .A2(new_n457_), .A3(new_n453_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .A4(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n557_), .A2(new_n725_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n572_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n735_), .B1(new_n747_), .B2(KEYINPUT57), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n740_), .A2(new_n741_), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n737_), .A2(new_n738_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n749_), .A2(new_n750_), .B1(new_n557_), .B2(new_n725_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n572_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n482_), .B1(new_n748_), .B2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n535_), .A2(new_n562_), .A3(new_n458_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n535_), .A2(new_n562_), .A3(new_n458_), .A4(new_n756_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n754_), .A2(new_n761_), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n313_), .B(new_n593_), .C1(new_n397_), .C2(new_n396_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT59), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n748_), .A2(KEYINPUT120), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n747_), .A2(KEYINPUT57), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT120), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n735_), .C1(new_n747_), .C2(KEYINPUT57), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n482_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n761_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n763_), .A2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n763_), .A2(new_n774_), .ZN(new_n776_));
  OR3_X1    g575(.A1(new_n775_), .A2(new_n776_), .A3(KEYINPUT59), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n765_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G113gat), .B1(new_n778_), .B2(new_n458_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n458_), .A2(G113gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n764_), .B2(new_n780_), .ZN(G1340gat));
  OAI21_X1  g580(.A(G120gat), .B1(new_n778_), .B2(new_n562_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT60), .ZN(new_n783_));
  AOI21_X1  g582(.A(G120gat), .B1(new_n563_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT121), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n783_), .B2(G120gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n785_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n782_), .B1(new_n764_), .B2(new_n788_), .ZN(G1341gat));
  OAI21_X1  g588(.A(G127gat), .B1(new_n778_), .B2(new_n482_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n482_), .A2(G127gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n764_), .B2(new_n791_), .ZN(G1342gat));
  OAI21_X1  g591(.A(G134gat), .B1(new_n778_), .B2(new_n615_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n573_), .A2(G134gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n764_), .B2(new_n794_), .ZN(G1343gat));
  NOR4_X1   g594(.A1(new_n399_), .A2(new_n582_), .A3(new_n387_), .A4(new_n313_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n762_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n459_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n563_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g601(.A1(new_n797_), .A2(new_n482_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT61), .B(G155gat), .Z(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(G1346gat));
  OR3_X1    g604(.A1(new_n797_), .A2(G162gat), .A3(new_n573_), .ZN(new_n806_));
  OAI21_X1  g605(.A(G162gat), .B1(new_n797_), .B2(new_n615_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1347gat));
  NOR2_X1   g607(.A1(new_n583_), .A2(new_n314_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n420_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n753_), .B1(new_n748_), .B2(KEYINPUT120), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n481_), .B1(new_n812_), .B2(new_n769_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n459_), .B(new_n811_), .C1(new_n813_), .C2(new_n760_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT122), .B1(new_n814_), .B2(G169gat), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT62), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n772_), .A2(new_n811_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n459_), .A2(new_n336_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT123), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n815_), .A2(new_n816_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n815_), .A2(new_n816_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n814_), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(G1348gat));
  NAND3_X1  g622(.A1(new_n772_), .A2(new_n563_), .A3(new_n811_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n230_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT124), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n752_), .B1(new_n751_), .B2(new_n572_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n767_), .A3(new_n735_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n760_), .B1(new_n828_), .B2(new_n482_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n826_), .B1(new_n829_), .B2(new_n420_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n762_), .A2(KEYINPUT124), .A3(new_n387_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n562_), .A2(new_n212_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n809_), .A4(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n825_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT125), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n825_), .A2(new_n833_), .A3(KEYINPUT125), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1349gat));
  NAND4_X1  g637(.A1(new_n830_), .A2(new_n831_), .A3(new_n481_), .A4(new_n809_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(new_n206_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n481_), .A2(new_n333_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n811_), .B(new_n841_), .C1(new_n813_), .C2(new_n760_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT126), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n772_), .A2(KEYINPUT126), .A3(new_n811_), .A4(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT127), .B1(new_n840_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(new_n206_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT127), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(G1350gat));
  NAND4_X1  g650(.A1(new_n817_), .A2(new_n203_), .A3(new_n205_), .A4(new_n572_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n817_), .A2(new_n616_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n202_), .ZN(G1351gat));
  NOR4_X1   g653(.A1(new_n583_), .A2(new_n399_), .A3(new_n387_), .A4(new_n567_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n762_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n459_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n563_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n481_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n863_));
  AND2_X1   g662(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n862_), .B2(new_n863_), .ZN(G1354gat));
  OR3_X1    g665(.A1(new_n856_), .A2(G218gat), .A3(new_n573_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G218gat), .B1(new_n856_), .B2(new_n615_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1355gat));
endmodule


