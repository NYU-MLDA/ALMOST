//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  OAI21_X1  g000(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(new_n202_), .B1(G169gat), .B2(G176gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT82), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(KEYINPUT82), .ZN(new_n205_));
  NOR3_X1   g004(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n205_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT83), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n214_), .B2(new_n211_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n217_), .A2(KEYINPUT85), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(KEYINPUT85), .ZN(new_n219_));
  OAI21_X1  g018(.A(G169gat), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT86), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT22), .B1(KEYINPUT84), .B2(G169gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(KEYINPUT84), .B2(G169gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT86), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n225_), .B(G169gat), .C1(new_n218_), .C2(new_n219_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT87), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n230_), .B1(new_n214_), .B2(KEYINPUT23), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(G183gat), .B2(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT87), .B1(new_n227_), .B2(new_n228_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n216_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G99gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n235_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G113gat), .B(G120gat), .Z(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n238_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(G15gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT30), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT31), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n243_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n243_), .A2(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT93), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT21), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n256_), .ZN(new_n260_));
  MUX2_X1   g059(.A(new_n257_), .B(new_n260_), .S(new_n254_), .Z(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(KEYINPUT21), .B2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G141gat), .B(G148gat), .Z(new_n263_));
  AND3_X1   g062(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT1), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n267_));
  OR2_X1    g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n264_), .A2(new_n265_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(KEYINPUT1), .B2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n267_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n263_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n270_), .A2(new_n268_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT2), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT3), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT3), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n275_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n276_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n276_), .A2(new_n284_), .ZN(new_n286_));
  AND4_X1   g085(.A1(new_n275_), .A2(new_n285_), .A3(new_n282_), .A4(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n274_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n273_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n253_), .B(new_n262_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n273_), .B2(new_n288_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n261_), .A2(KEYINPUT21), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(KEYINPUT21), .B2(new_n258_), .ZN(new_n294_));
  OAI211_X1 g093(.A(G228gat), .B(G233gat), .C1(new_n292_), .C2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G78gat), .B(G106gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n300_), .A2(KEYINPUT94), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G22gat), .B(G50gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT92), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n273_), .A2(new_n288_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n308_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n305_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n289_), .A2(new_n306_), .A3(new_n290_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT28), .B1(new_n308_), .B2(KEYINPUT29), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(new_n304_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n301_), .B1(new_n302_), .B2(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n310_), .A2(new_n313_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT94), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n300_), .A4(new_n298_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n252_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT99), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n273_), .A2(new_n288_), .A3(new_n242_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n242_), .B1(new_n273_), .B2(new_n288_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n308_), .A2(new_n325_), .A3(new_n241_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n322_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n324_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n273_), .A2(new_n288_), .A3(new_n242_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n328_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(KEYINPUT4), .A3(new_n333_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n328_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT99), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n331_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G57gat), .B(G85gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT101), .ZN(new_n340_));
  INV_X1    g139(.A(G1gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n343_));
  INV_X1    g142(.A(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n342_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n346_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n331_), .A2(new_n337_), .A3(new_n348_), .A4(new_n334_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT20), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G169gat), .ZN(new_n353_));
  INV_X1    g152(.A(G176gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n228_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(KEYINPUT96), .A3(new_n228_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n358_), .B(new_n359_), .C1(new_n215_), .C2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n203_), .A2(new_n206_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n208_), .B(KEYINPUT95), .ZN(new_n363_));
  INV_X1    g162(.A(new_n207_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n231_), .B(new_n362_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT103), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n262_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n361_), .A2(KEYINPUT103), .A3(new_n365_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n352_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n235_), .A2(new_n262_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT19), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n294_), .B(new_n216_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n352_), .B1(new_n366_), .B2(new_n262_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(new_n374_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT98), .ZN(new_n383_));
  XOR2_X1   g182(.A(G8gat), .B(G36gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n387_), .B(KEYINPUT104), .Z(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n378_), .A2(new_n374_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n371_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n374_), .ZN(new_n392_));
  OAI211_X1 g191(.A(KEYINPUT20), .B(new_n392_), .C1(new_n366_), .C2(new_n262_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n390_), .B(new_n387_), .C1(new_n391_), .C2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(KEYINPUT27), .ZN(new_n395_));
  INV_X1    g194(.A(new_n387_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n393_), .B1(new_n235_), .B2(new_n262_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n392_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT105), .B(KEYINPUT27), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n389_), .A2(new_n395_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n321_), .A2(new_n351_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT102), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n349_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n346_), .A2(new_n406_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n331_), .A2(new_n337_), .A3(new_n334_), .A4(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n335_), .A2(new_n328_), .A3(new_n327_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n332_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n346_), .A3(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n409_), .A2(new_n394_), .A3(new_n399_), .A4(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n405_), .B1(new_n407_), .B2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n394_), .A2(new_n412_), .A3(new_n399_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n349_), .A2(new_n406_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n415_), .A2(KEYINPUT102), .A3(new_n416_), .A4(new_n409_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n387_), .A2(KEYINPUT32), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n418_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n381_), .B2(new_n418_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n350_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n414_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n319_), .A2(new_n350_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n422_), .A2(new_n319_), .B1(new_n423_), .B2(new_n403_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n252_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n404_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G29gat), .B(G36gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT73), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G43gat), .B(G50gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n427_), .A2(KEYINPUT73), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(KEYINPUT73), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n429_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G15gat), .B(G22gat), .ZN(new_n437_));
  INV_X1    g236(.A(G8gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(new_n341_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G1gat), .B(G8gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G229gat), .A2(G233gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT15), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n435_), .B(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n442_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n435_), .B(new_n442_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n445_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G113gat), .B(G141gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G169gat), .B(G197gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  OR2_X1    g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n456_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n459_), .B(KEYINPUT81), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n426_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G232gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT34), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT6), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(G99gat), .A3(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT69), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  INV_X1    g274(.A(G99gat), .ZN(new_n476_));
  INV_X1    g275(.A(G106gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n473_), .A2(new_n474_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G85gat), .ZN(new_n482_));
  INV_X1    g281(.A(G92gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n484_), .A2(KEYINPUT67), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT67), .B1(new_n484_), .B2(new_n485_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT8), .B1(new_n481_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n470_), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n468_), .A2(KEYINPUT6), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n469_), .A2(new_n471_), .A3(KEYINPUT66), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n480_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n490_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n469_), .A2(new_n471_), .A3(KEYINPUT66), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT66), .B1(new_n469_), .B2(new_n471_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n478_), .B(new_n479_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n484_), .A2(new_n485_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n484_), .A2(KEYINPUT67), .A3(new_n485_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT8), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(new_n507_), .A3(KEYINPUT68), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n489_), .A2(new_n499_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT70), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT10), .B(G99gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT64), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n477_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n494_), .A2(new_n495_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT65), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n484_), .A2(new_n515_), .A3(KEYINPUT9), .ZN(new_n516_));
  OAI211_X1 g315(.A(G85gat), .B(G92gat), .C1(new_n515_), .C2(KEYINPUT9), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n509_), .A2(new_n510_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n510_), .B1(new_n509_), .B2(new_n519_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n435_), .B(KEYINPUT15), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n509_), .A2(new_n519_), .ZN(new_n524_));
  OAI22_X1  g323(.A1(new_n524_), .A2(new_n435_), .B1(KEYINPUT35), .B2(new_n464_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n467_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(KEYINPUT70), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n509_), .A2(new_n510_), .A3(new_n519_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n448_), .A3(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n509_), .A2(new_n519_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n530_), .A2(new_n436_), .B1(new_n466_), .B2(new_n465_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n467_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G134gat), .B(G162gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(KEYINPUT36), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n526_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n536_), .B(KEYINPUT36), .Z(new_n541_));
  AND3_X1   g340(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n532_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(new_n539_), .A3(new_n538_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT75), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n549_), .B2(KEYINPUT37), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT37), .ZN(new_n551_));
  AOI211_X1 g350(.A(KEYINPUT76), .B(new_n551_), .C1(new_n544_), .C2(new_n548_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n546_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n541_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n526_), .B2(new_n533_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT37), .B1(new_n555_), .B2(KEYINPUT75), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT76), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n547_), .B(KEYINPUT37), .C1(new_n555_), .C2(KEYINPUT75), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n557_), .A2(new_n545_), .A3(new_n540_), .A4(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n562_));
  XOR2_X1   g361(.A(G71gat), .B(G78gat), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT12), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n567_), .B2(new_n566_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n527_), .A2(new_n528_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n509_), .A2(new_n566_), .A3(new_n519_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT12), .ZN(new_n572_));
  INV_X1    g371(.A(new_n566_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n524_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n571_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G120gat), .B(G148gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n586_), .B(new_n587_), .C1(KEYINPUT72), .C2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT17), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n442_), .B(new_n602_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(new_n573_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n573_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT79), .ZN(new_n607_));
  AOI211_X1 g406(.A(new_n600_), .B(new_n601_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n604_), .A2(KEYINPUT79), .A3(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(KEYINPUT71), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n567_), .A3(new_n605_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n600_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT78), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n610_), .A2(KEYINPUT78), .A3(new_n600_), .A4(new_n611_), .ZN(new_n615_));
  AOI221_X4 g414(.A(KEYINPUT80), .B1(new_n608_), .B2(new_n609_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT80), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n609_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n553_), .A2(new_n559_), .A3(new_n593_), .A4(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n462_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT106), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n351_), .A2(KEYINPUT107), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n351_), .A2(KEYINPUT107), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n341_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n546_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n426_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n593_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n459_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n618_), .A2(new_n619_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n635_), .A2(new_n636_), .A3(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n634_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G1gat), .B1(new_n641_), .B2(new_n351_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n630_), .A2(new_n631_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n632_), .A2(new_n642_), .A3(new_n643_), .ZN(G1324gat));
  INV_X1    g443(.A(new_n403_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n625_), .A2(new_n438_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n640_), .A2(new_n645_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(G8gat), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT39), .B(new_n438_), .C1(new_n640_), .C2(new_n645_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n646_), .B(new_n652_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  AOI21_X1  g455(.A(new_n245_), .B1(new_n640_), .B2(new_n425_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT41), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n625_), .A2(new_n245_), .A3(new_n425_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1326gat));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n640_), .B2(new_n320_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT42), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n625_), .A2(new_n661_), .A3(new_n320_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1327gat));
  NOR3_X1   g464(.A1(new_n635_), .A2(new_n621_), .A3(new_n633_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n462_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G29gat), .B1(new_n667_), .B2(new_n350_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n635_), .A2(new_n636_), .A3(new_n621_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n553_), .A2(new_n559_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n426_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n426_), .B2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(KEYINPUT44), .B(new_n669_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n628_), .A2(new_n344_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n668_), .B1(new_n678_), .B2(new_n679_), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n676_), .A2(new_n645_), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  NOR2_X1   g481(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n403_), .A2(G36gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n462_), .A2(new_n666_), .A3(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT45), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n682_), .A2(new_n684_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT110), .Z(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n682_), .A2(new_n690_), .A3(new_n684_), .A4(new_n687_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1329gat));
  INV_X1    g493(.A(G43gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n252_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n676_), .A2(new_n677_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT111), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n676_), .A2(new_n699_), .A3(new_n677_), .A4(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n667_), .A2(new_n425_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n695_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT47), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n698_), .A2(new_n705_), .A3(new_n700_), .A4(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1330gat));
  INV_X1    g506(.A(G50gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n667_), .A2(new_n708_), .A3(new_n320_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n676_), .A2(new_n320_), .A3(new_n677_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n710_), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT112), .B1(new_n710_), .B2(G50gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1331gat));
  INV_X1    g512(.A(new_n621_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n461_), .A2(new_n714_), .A3(new_n593_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n634_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n351_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n426_), .A2(new_n636_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n671_), .ZN(new_n720_));
  AND4_X1   g519(.A1(new_n635_), .A2(new_n719_), .A3(new_n621_), .A4(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n629_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n716_), .B2(new_n645_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT48), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n721_), .A2(new_n725_), .A3(new_n645_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n716_), .B2(new_n425_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT49), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n721_), .A2(new_n730_), .A3(new_n425_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1334gat));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n716_), .B2(new_n320_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT50), .Z(new_n737_));
  NAND3_X1  g536(.A1(new_n721_), .A2(new_n735_), .A3(new_n320_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1335gat));
  NAND2_X1  g538(.A1(new_n635_), .A2(new_n714_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n633_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n719_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n482_), .A3(new_n629_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n672_), .A2(new_n673_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(new_n459_), .A3(new_n740_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n350_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n747_), .B2(new_n482_), .ZN(G1336gat));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n483_), .A3(new_n645_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n745_), .A2(new_n645_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n751_), .B2(new_n483_), .ZN(G1337gat));
  XNOR2_X1  g551(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n742_), .A2(new_n425_), .A3(new_n512_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n476_), .B1(new_n745_), .B2(new_n425_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n755_), .B(KEYINPUT113), .ZN(new_n760_));
  INV_X1    g559(.A(new_n758_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n753_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1338gat));
  NAND4_X1  g562(.A1(new_n719_), .A2(new_n477_), .A3(new_n320_), .A4(new_n741_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT115), .Z(new_n765_));
  NOR2_X1   g564(.A1(new_n740_), .A2(new_n459_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n320_), .B(new_n766_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n767_), .A2(G106gat), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n767_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n765_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n765_), .B(new_n774_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT124), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n444_), .B(new_n451_), .C1(new_n522_), .C2(new_n443_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n456_), .B1(new_n450_), .B2(new_n445_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n453_), .A2(new_n456_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n586_), .A2(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT122), .Z(new_n782_));
  NOR2_X1   g581(.A1(new_n576_), .A2(KEYINPUT120), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n570_), .A2(new_n575_), .A3(new_n783_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n579_), .A2(KEYINPUT55), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n570_), .A2(new_n575_), .A3(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n786_), .B2(new_n783_), .ZN(new_n787_));
  XOR2_X1   g586(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n788_));
  NAND2_X1  g587(.A1(new_n577_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT119), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n577_), .A2(new_n791_), .A3(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n585_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n782_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n782_), .A2(new_n798_), .A3(KEYINPUT58), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n671_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n586_), .A2(new_n459_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n797_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n585_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n588_), .A2(new_n780_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n546_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n810_), .A2(KEYINPUT121), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n804_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n809_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n633_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT57), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n803_), .B1(new_n812_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n623_), .B2(new_n460_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  NOR4_X1   g620(.A1(new_n622_), .A2(new_n821_), .A3(KEYINPUT54), .A4(new_n461_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n622_), .A2(new_n461_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n819_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n821_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n818_), .A2(new_n714_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n628_), .A2(new_n645_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n321_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT123), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n829_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n777_), .B1(new_n827_), .B2(new_n835_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n818_), .A2(new_n638_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT59), .B1(new_n837_), .B2(new_n829_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n835_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(new_n824_), .B2(new_n819_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n840_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n811_), .B1(new_n810_), .B2(KEYINPUT121), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n815_), .A2(new_n816_), .A3(KEYINPUT57), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n621_), .B1(new_n844_), .B2(new_n803_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n839_), .B(KEYINPUT124), .C1(new_n841_), .C2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n836_), .A2(new_n838_), .A3(new_n461_), .A4(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G113gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n841_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n818_), .A2(new_n638_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n830_), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n852_), .A2(G113gat), .A3(new_n636_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n848_), .A2(new_n853_), .ZN(G1340gat));
  NAND4_X1  g653(.A1(new_n836_), .A2(new_n838_), .A3(new_n635_), .A4(new_n846_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G120gat), .ZN(new_n856_));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(KEYINPUT60), .B2(new_n857_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n852_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n860_), .ZN(G1341gat));
  NAND4_X1  g660(.A1(new_n836_), .A2(new_n838_), .A3(new_n637_), .A4(new_n846_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G127gat), .ZN(new_n863_));
  OR3_X1    g662(.A1(new_n852_), .A2(G127gat), .A3(new_n714_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1342gat));
  XOR2_X1   g664(.A(KEYINPUT125), .B(G134gat), .Z(new_n866_));
  NOR2_X1   g665(.A1(new_n720_), .A2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n836_), .A2(new_n838_), .A3(new_n846_), .A4(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(G134gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n852_), .B2(new_n633_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1343gat));
  NOR2_X1   g670(.A1(new_n425_), .A2(new_n319_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n851_), .A2(new_n459_), .A3(new_n828_), .A4(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g673(.A1(new_n851_), .A2(new_n635_), .A3(new_n828_), .A4(new_n872_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g675(.A1(new_n851_), .A2(new_n621_), .A3(new_n828_), .A4(new_n872_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  NOR3_X1   g678(.A1(new_n837_), .A2(new_n425_), .A3(new_n319_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n880_), .A2(new_n828_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n671_), .A2(G162gat), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT126), .Z(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n546_), .A3(new_n828_), .ZN(new_n884_));
  INV_X1    g683(.A(G162gat), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n881_), .A2(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n252_), .A2(new_n403_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n628_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n320_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n459_), .B(new_n889_), .C1(new_n845_), .C2(new_n841_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n890_), .A2(new_n891_), .A3(G169gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n890_), .B2(G169gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n889_), .B1(new_n845_), .B2(new_n841_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n459_), .A2(new_n353_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT127), .ZN(new_n896_));
  OAI22_X1  g695(.A1(new_n892_), .A2(new_n893_), .B1(new_n894_), .B2(new_n896_), .ZN(G1348gat));
  INV_X1    g696(.A(new_n894_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G176gat), .B1(new_n898_), .B2(new_n635_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n837_), .A2(new_n320_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n888_), .A2(new_n354_), .A3(new_n593_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  NOR3_X1   g701(.A1(new_n894_), .A2(new_n207_), .A3(new_n638_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n900_), .A2(new_n621_), .A3(new_n628_), .A4(new_n887_), .ZN(new_n904_));
  INV_X1    g703(.A(G183gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n894_), .B2(new_n720_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n633_), .A2(new_n363_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n894_), .B2(new_n908_), .ZN(G1351gat));
  NOR2_X1   g708(.A1(new_n403_), .A2(new_n350_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n851_), .A2(new_n459_), .A3(new_n872_), .A4(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g711(.A1(new_n851_), .A2(new_n635_), .A3(new_n872_), .A4(new_n910_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g713(.A1(new_n851_), .A2(new_n637_), .A3(new_n872_), .A4(new_n910_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT63), .B(G211gat), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n915_), .B2(new_n918_), .ZN(G1354gat));
  NAND4_X1  g718(.A1(new_n851_), .A2(new_n671_), .A3(new_n872_), .A4(new_n910_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G218gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n880_), .A2(new_n910_), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n633_), .A2(G218gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1355gat));
endmodule


