//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT10), .B(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  OR3_X1    g006(.A1(new_n206_), .A2(new_n207_), .A3(G106gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT66), .A3(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n211_), .A2(new_n213_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n209_), .A2(KEYINPUT66), .A3(KEYINPUT9), .A4(new_n210_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n207_), .B1(new_n206_), .B2(G106gat), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n208_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223_));
  OAI22_X1  g022(.A1(new_n223_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .A4(KEYINPUT67), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n216_), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n224_), .B(new_n228_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n232_));
  AND2_X1   g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n232_), .B1(new_n233_), .B2(new_n212_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n209_), .A2(KEYINPUT68), .A3(new_n210_), .ZN(new_n235_));
  AND4_X1   g034(.A1(new_n222_), .A2(new_n231_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n235_), .A2(new_n234_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n222_), .B1(new_n237_), .B2(new_n231_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n221_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n205_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G232gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT34), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(KEYINPUT69), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n244_), .B(new_n221_), .C1(new_n236_), .C2(new_n238_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n204_), .ZN(new_n247_));
  OAI221_X1 g046(.A(new_n240_), .B1(KEYINPUT35), .B2(new_n242_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n242_), .A2(KEYINPUT35), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G190gat), .B(G218gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G134gat), .B(G162gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT36), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n253_), .A2(KEYINPUT36), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT37), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT71), .B(G15gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(G22gat), .ZN(new_n262_));
  INV_X1    g061(.A(G1gat), .ZN(new_n263_));
  INV_X1    g062(.A(G8gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT14), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G8gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G57gat), .B(G64gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G71gat), .B(G78gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT11), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(new_n272_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n273_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n270_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT74), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G127gat), .B(G155gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G183gat), .B(G211gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT17), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n285_), .A2(new_n287_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n279_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n279_), .A2(new_n288_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT75), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n260_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G113gat), .B(G141gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G169gat), .B(G197gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n268_), .A2(new_n205_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT76), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n268_), .A2(new_n247_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G229gat), .A2(G233gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n268_), .B(new_n247_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n297_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n297_), .ZN(new_n310_));
  AOI211_X1 g109(.A(KEYINPUT77), .B(new_n310_), .C1(new_n304_), .C2(new_n306_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT25), .B(G183gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT26), .B(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT24), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(G169gat), .B2(G176gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT24), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT78), .B1(new_n324_), .B2(new_n320_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n316_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT79), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n316_), .A2(new_n322_), .A3(new_n325_), .A4(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(new_n317_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n330_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n327_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT80), .B(G176gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT22), .B(G169gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n333_), .B(new_n334_), .C1(G183gat), .C2(G190gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n323_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G71gat), .B(G99gat), .ZN(new_n343_));
  INV_X1    g142(.A(G43gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n342_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(G15gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT30), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT83), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n335_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n326_), .B2(KEYINPUT79), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n337_), .A2(new_n338_), .B1(G169gat), .B2(G176gat), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n355_), .A2(new_n329_), .B1(new_n340_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(new_n345_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n351_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G113gat), .B(G120gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G134gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G127gat), .ZN(new_n364_));
  INV_X1    g163(.A(G127gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G134gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n362_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n365_), .A2(G134gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n363_), .A2(G127gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n361_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT31), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n360_), .A2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n353_), .B(new_n359_), .C1(new_n378_), .C2(new_n377_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT84), .Z(new_n385_));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT19), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT20), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n314_), .A2(new_n315_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n335_), .A2(new_n395_), .B1(new_n356_), .B2(new_n340_), .ZN(new_n396_));
  INV_X1    g195(.A(G197gat), .ZN(new_n397_));
  INV_X1    g196(.A(G204gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G197gat), .A2(G204gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(KEYINPUT21), .A3(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G211gat), .B(G218gat), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT21), .ZN(new_n404_));
  INV_X1    g203(.A(new_n400_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G197gat), .A2(G204gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n394_), .B1(new_n396_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n357_), .B2(new_n409_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT20), .B1(new_n396_), .B2(new_n409_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n357_), .B2(new_n409_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n391_), .B(new_n411_), .C1(new_n413_), .C2(new_n393_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT93), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT92), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n390_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n403_), .A2(new_n408_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n395_), .A2(new_n335_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n341_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n421_), .B2(KEYINPUT90), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n396_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n418_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n342_), .A2(new_n419_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n393_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n336_), .A2(new_n341_), .A3(new_n409_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n418_), .B1(new_n421_), .B2(new_n419_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n428_), .A2(new_n393_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n417_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n429_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n393_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n391_), .A4(new_n411_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n415_), .A2(new_n431_), .A3(KEYINPUT27), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT27), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n391_), .B1(new_n434_), .B2(new_n411_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n393_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT20), .B(new_n393_), .C1(new_n421_), .C2(new_n419_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n342_), .B2(new_n419_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n440_), .A2(new_n442_), .A3(new_n390_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n438_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G141gat), .A2(G148gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G141gat), .A2(G148gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT2), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n447_), .A2(new_n450_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G155gat), .A2(G162gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n448_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(new_n445_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT85), .B1(new_n456_), .B2(KEYINPUT1), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n456_), .A2(KEYINPUT1), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n454_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n458_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT28), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT29), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n463_), .A2(new_n454_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n462_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n465_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n460_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n457_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT28), .B1(new_n475_), .B2(KEYINPUT29), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n470_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT86), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n409_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT87), .B(KEYINPUT29), .Z(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n467_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n469_), .B1(new_n474_), .B2(new_n457_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n484_), .B1(new_n488_), .B2(new_n409_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G22gat), .B(G50gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n482_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n494_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n496_), .A2(new_n481_), .A3(new_n479_), .A4(new_n492_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n376_), .B1(new_n458_), .B2(new_n466_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n474_), .A2(new_n375_), .A3(new_n370_), .A4(new_n457_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT4), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT4), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n475_), .A2(new_n504_), .A3(new_n376_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n499_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G1gat), .B(G29gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G85gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT0), .B(G57gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n499_), .A2(KEYINPUT4), .A3(new_n500_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n505_), .A2(new_n503_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n507_), .B(new_n514_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n437_), .A2(new_n444_), .A3(new_n498_), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT94), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n497_), .B2(new_n495_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n444_), .A4(new_n437_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT89), .B1(new_n439_), .B2(new_n443_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n499_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n512_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n505_), .A2(new_n502_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n501_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n517_), .A2(KEYINPUT33), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT33), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n506_), .A2(new_n531_), .A3(new_n507_), .A4(new_n514_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n529_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n390_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n414_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n525_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n391_), .A2(KEYINPUT32), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n434_), .A2(new_n411_), .A3(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n427_), .A2(new_n430_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n518_), .B(new_n539_), .C1(new_n540_), .C2(new_n538_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n498_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n521_), .B(new_n524_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n385_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n384_), .B(KEYINPUT84), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n437_), .A2(new_n444_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(new_n498_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n519_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n313_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n243_), .A2(new_n245_), .A3(new_n277_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n278_), .A2(KEYINPUT12), .A3(new_n239_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT64), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n245_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n215_), .A2(new_n217_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n559_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n235_), .A2(new_n234_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT8), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n237_), .A2(new_n222_), .A3(new_n231_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n244_), .B1(new_n564_), .B2(new_n221_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n278_), .B1(new_n558_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n554_), .A2(new_n557_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n552_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n556_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n569_), .A2(new_n571_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(KEYINPUT70), .A3(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT13), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n582_), .A2(KEYINPUT13), .A3(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n294_), .A2(new_n551_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT95), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n263_), .A3(new_n518_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT38), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n292_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n312_), .A3(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT96), .ZN(new_n597_));
  INV_X1    g396(.A(new_n258_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(KEYINPUT96), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n519_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n592_), .A2(new_n593_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(new_n602_), .A3(new_n603_), .ZN(G1324gat));
  XNOR2_X1  g403(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n605_));
  INV_X1    g404(.A(new_n548_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n607_), .A2(new_n608_), .A3(G8gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n607_), .B2(G8gat), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n591_), .A2(new_n264_), .A3(new_n548_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n605_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n612_), .B(new_n605_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(G1325gat));
  INV_X1    g415(.A(KEYINPUT41), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n601_), .A2(new_n385_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(G15gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n618_), .B2(G15gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n617_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(G15gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT98), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(KEYINPUT41), .A3(new_n620_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n591_), .A2(new_n348_), .A3(new_n547_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT99), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n623_), .A2(new_n626_), .A3(new_n630_), .A4(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(G1326gat));
  INV_X1    g431(.A(new_n498_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G22gat), .B1(new_n601_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(G22gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT100), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n591_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n293_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n640_), .A2(new_n588_), .A3(new_n258_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n551_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n642_), .A2(G29gat), .A3(new_n519_), .ZN(new_n643_));
  XOR2_X1   g442(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n546_), .A2(new_n550_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n260_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n645_), .A2(KEYINPUT101), .A3(new_n646_), .A4(new_n260_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(new_n260_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT43), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n649_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n640_), .A2(new_n588_), .A3(new_n313_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n644_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT104), .B(new_n644_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n655_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n519_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n662_), .A2(KEYINPUT105), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT105), .B1(new_n662_), .B2(new_n665_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n643_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  NOR3_X1   g468(.A1(new_n642_), .A2(G36gat), .A3(new_n606_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n663_), .A2(new_n548_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n674_));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT46), .B(new_n672_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1329gat));
  NOR2_X1   g479(.A1(new_n385_), .A2(new_n344_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n664_), .B(new_n682_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n641_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT107), .B(G43gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT47), .B1(new_n683_), .B2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n664_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n681_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n686_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(G1330gat));
  INV_X1    g492(.A(G50gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n633_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n641_), .A2(new_n498_), .A3(new_n551_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n689_), .A2(new_n695_), .B1(new_n694_), .B2(new_n696_), .ZN(G1331gat));
  NAND4_X1  g496(.A1(new_n599_), .A2(new_n313_), .A3(new_n588_), .A4(new_n640_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n519_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n312_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n294_), .A2(new_n700_), .A3(new_n588_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n519_), .A2(G57gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(G1332gat));
  OAI21_X1  g502(.A(G64gat), .B1(new_n698_), .B2(new_n606_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT48), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n606_), .A2(G64gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n701_), .B2(new_n706_), .ZN(G1333gat));
  OAI21_X1  g506(.A(G71gat), .B1(new_n698_), .B2(new_n385_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n385_), .A2(G71gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n701_), .B2(new_n711_), .ZN(G1334gat));
  OAI21_X1  g511(.A(G78gat), .B1(new_n698_), .B2(new_n633_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT50), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n633_), .A2(G78gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n701_), .B2(new_n715_), .ZN(G1335gat));
  AND4_X1   g515(.A1(new_n588_), .A2(new_n700_), .A3(new_n293_), .A4(new_n598_), .ZN(new_n717_));
  INV_X1    g516(.A(G85gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n518_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n589_), .A2(new_n640_), .A3(new_n312_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n653_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT109), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(new_n518_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n723_), .B2(new_n718_), .ZN(G1336gat));
  AOI21_X1  g523(.A(G92gat), .B1(new_n717_), .B2(new_n548_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n548_), .A2(G92gat), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT110), .Z(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n722_), .B2(new_n727_), .ZN(G1337gat));
  NAND3_X1  g527(.A1(new_n653_), .A2(new_n547_), .A3(new_n720_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n385_), .A2(new_n206_), .ZN(new_n730_));
  AOI22_X1  g529(.A1(new_n729_), .A2(G99gat), .B1(new_n717_), .B2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(G1338gat));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n653_), .A2(new_n498_), .A3(new_n720_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT113), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n653_), .A2(new_n738_), .A3(new_n498_), .A4(new_n720_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G106gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n734_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n736_), .A2(KEYINPUT114), .A3(G106gat), .A4(new_n739_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(KEYINPUT52), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n734_), .B(new_n744_), .C1(new_n737_), .C2(new_n740_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n717_), .A2(new_n227_), .A3(new_n498_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT112), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n743_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT53), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n743_), .A2(new_n750_), .A3(new_n745_), .A4(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1339gat));
  NAND3_X1  g551(.A1(new_n547_), .A2(new_n518_), .A3(new_n549_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n312_), .A2(new_n579_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n554_), .A2(new_n755_), .A3(new_n568_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT12), .B1(new_n246_), .B2(new_n278_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n552_), .A2(new_n553_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT116), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n759_), .A3(new_n556_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT117), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n277_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n552_), .B(new_n553_), .C1(new_n763_), .C2(KEYINPUT12), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(new_n556_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n554_), .A2(new_n568_), .A3(KEYINPUT55), .A4(new_n557_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n756_), .A2(new_n759_), .A3(new_n768_), .A4(new_n556_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n761_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n576_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(KEYINPUT56), .A3(new_n576_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n754_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n299_), .B(new_n302_), .C1(new_n268_), .C2(new_n247_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n305_), .A2(new_n301_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n297_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n307_), .B2(new_n297_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT57), .B(new_n258_), .C1(new_n775_), .C2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT118), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n258_), .B1(new_n775_), .B2(new_n780_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n774_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n770_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n576_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n773_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(new_n579_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n779_), .A2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n790_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n791_), .B1(new_n790_), .B2(new_n793_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT120), .B(new_n260_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n783_), .A2(KEYINPUT118), .A3(new_n784_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n786_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n795_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n790_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT120), .B1(new_n801_), .B2(new_n260_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n292_), .B1(new_n798_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n294_), .A2(new_n313_), .A3(new_n589_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n753_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n312_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  INV_X1    g609(.A(new_n753_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n812_), .B2(new_n811_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n806_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n801_), .A2(new_n260_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n785_), .A2(new_n781_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n640_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n814_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n807_), .B2(new_n810_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT122), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT122), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n819_), .C1(new_n807_), .C2(new_n810_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n313_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n809_), .B1(new_n824_), .B2(new_n808_), .ZN(G1340gat));
  XOR2_X1   g624(.A(KEYINPUT123), .B(G120gat), .Z(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n589_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n753_), .B(new_n828_), .C1(new_n803_), .C2(new_n806_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT124), .Z(new_n830_));
  INV_X1    g629(.A(new_n826_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n820_), .B2(new_n589_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n807_), .B2(new_n640_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n821_), .A2(new_n823_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT125), .B(G127gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n292_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n834_), .B1(new_n835_), .B2(new_n837_), .ZN(G1342gat));
  NAND3_X1  g637(.A1(new_n807_), .A2(new_n363_), .A3(new_n598_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n260_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n841_), .B2(new_n363_), .ZN(G1343gat));
  AOI21_X1  g641(.A(new_n547_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(new_n518_), .A3(new_n606_), .A4(new_n498_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n313_), .ZN(new_n845_));
  INV_X1    g644(.A(G141gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1344gat));
  NOR2_X1   g646(.A1(new_n844_), .A2(new_n589_), .ZN(new_n848_));
  INV_X1    g647(.A(G148gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1345gat));
  NOR2_X1   g649(.A1(new_n844_), .A2(new_n293_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT61), .B(G155gat), .Z(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  OAI21_X1  g652(.A(G162gat), .B1(new_n844_), .B2(new_n840_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n258_), .A2(G162gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n844_), .B2(new_n855_), .ZN(G1347gat));
  NOR2_X1   g655(.A1(new_n606_), .A2(new_n518_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n547_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n498_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n818_), .B2(new_n815_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT126), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n312_), .A3(new_n338_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n861_), .A2(new_n312_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(G169gat), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n868_), .A2(new_n867_), .A3(G169gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n866_), .B1(new_n869_), .B2(new_n870_), .ZN(G1348gat));
  NAND2_X1  g670(.A1(new_n865_), .A2(new_n588_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n498_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n873_));
  INV_X1    g672(.A(G176gat), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n589_), .A2(new_n874_), .A3(new_n858_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n872_), .A2(new_n337_), .B1(new_n873_), .B2(new_n875_), .ZN(G1349gat));
  NOR2_X1   g675(.A1(new_n292_), .A2(new_n314_), .ZN(new_n877_));
  INV_X1    g676(.A(G183gat), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n873_), .A2(new_n547_), .A3(new_n640_), .A4(new_n857_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n865_), .A2(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(G1350gat));
  NAND3_X1  g679(.A1(new_n865_), .A2(new_n315_), .A3(new_n598_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n840_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n882_));
  INV_X1    g681(.A(G190gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1351gat));
  NAND2_X1  g683(.A1(new_n548_), .A2(new_n522_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n843_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n313_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n397_), .ZN(G1352gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n589_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n398_), .ZN(G1353gat));
  OR2_X1    g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT63), .B(G211gat), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n887_), .A2(new_n292_), .ZN(new_n894_));
  MUX2_X1   g693(.A(new_n892_), .B(new_n893_), .S(new_n894_), .Z(G1354gat));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n887_), .A2(new_n896_), .A3(new_n840_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n887_), .A2(KEYINPUT127), .A3(new_n258_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(G218gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT127), .B1(new_n887_), .B2(new_n258_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n897_), .B1(new_n899_), .B2(new_n900_), .ZN(G1355gat));
endmodule


