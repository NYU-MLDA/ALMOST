//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  INV_X1    g000(.A(KEYINPUT107), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT10), .B(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT64), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(G106gat), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT9), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT9), .A3(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n213_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n209_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n206_), .A2(KEYINPUT64), .A3(new_n207_), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT64), .B1(new_n206_), .B2(new_n207_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n221_), .A2(new_n218_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n213_), .A4(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT7), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n234_), .B(new_n224_), .C1(new_n235_), .C2(KEYINPUT67), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(KEYINPUT67), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n218_), .A2(new_n233_), .A3(new_n236_), .A4(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n219_), .A2(new_n220_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n231_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n238_), .A2(new_n231_), .A3(new_n239_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n223_), .B(new_n230_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G64gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n244_));
  XOR2_X1   g043(.A(G71gat), .B(G78gat), .Z(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n242_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n242_), .A2(new_n249_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n252_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  AOI211_X1 g055(.A(KEYINPUT71), .B(new_n254_), .C1(new_n242_), .C2(new_n249_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n251_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n242_), .A2(KEYINPUT12), .A3(new_n249_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT69), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n260_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n250_), .B1(KEYINPUT68), .B2(new_n253_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(KEYINPUT68), .B2(new_n253_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n260_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G120gat), .B(G148gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(G176gat), .B(G204gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(new_n268_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT13), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(KEYINPUT13), .A3(new_n277_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G190gat), .B(G218gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT78), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G134gat), .B(G162gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT79), .B(KEYINPUT36), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT75), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G29gat), .B(G36gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n290_), .A2(KEYINPUT74), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(KEYINPUT74), .ZN(new_n292_));
  XOR2_X1   g091(.A(G43gat), .B(G50gat), .Z(new_n293_));
  OR3_X1    g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n289_), .B1(new_n242_), .B2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n223_), .A2(new_n230_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n241_), .A2(new_n240_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT75), .A4(new_n296_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT34), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(KEYINPUT35), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(KEYINPUT35), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT73), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT15), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n296_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT15), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n309_), .B1(new_n313_), .B2(new_n242_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n305_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n298_), .A2(new_n301_), .A3(KEYINPUT76), .A4(new_n304_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n242_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(KEYINPUT77), .A3(new_n309_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT77), .B1(new_n320_), .B2(new_n309_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n288_), .B(new_n315_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n309_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n327_), .A2(new_n321_), .B1(new_n306_), .B2(new_n314_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n286_), .B(KEYINPUT36), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n324_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT37), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G15gat), .B(G22gat), .ZN(new_n332_));
  INV_X1    g131(.A(G1gat), .ZN(new_n333_));
  INV_X1    g132(.A(G8gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT14), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G8gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(new_n249_), .Z(new_n339_));
  NAND2_X1  g138(.A1(G231gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G127gat), .B(G155gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT16), .ZN(new_n343_));
  XOR2_X1   g142(.A(G183gat), .B(G211gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT17), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n345_), .A2(new_n346_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n341_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n347_), .B2(new_n341_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT37), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n351_), .B(new_n324_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n282_), .A2(new_n331_), .A3(new_n350_), .A4(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n353_), .A2(KEYINPUT80), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(KEYINPUT80), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G127gat), .B(G134gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G113gat), .B(G120gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n356_), .A2(new_n357_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT89), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT31), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT88), .B(G15gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G183gat), .ZN(new_n369_));
  INV_X1    g168(.A(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT86), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT22), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(G169gat), .ZN(new_n377_));
  AOI21_X1  g176(.A(G176gat), .B1(new_n376_), .B2(G169gat), .ZN(new_n378_));
  INV_X1    g177(.A(G169gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n368_), .A2(new_n371_), .A3(new_n382_), .A4(new_n372_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n374_), .A2(new_n381_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  INV_X1    g185(.A(G176gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n379_), .A3(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n388_), .A2(new_n368_), .A3(new_n372_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT25), .B(G183gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT26), .B(G190gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n386_), .B1(G169gat), .B2(G176gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n379_), .A2(new_n387_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n390_), .A2(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n389_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n369_), .A2(KEYINPUT25), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT25), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G183gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n370_), .A2(KEYINPUT26), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT26), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G190gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .A4(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n393_), .A2(KEYINPUT24), .A3(new_n384_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n395_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT87), .B(new_n385_), .C1(new_n396_), .C2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT84), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n405_), .A3(new_n389_), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT87), .B1(new_n411_), .B2(new_n385_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n365_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414_));
  INV_X1    g213(.A(G43gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n385_), .B1(new_n396_), .B2(new_n406_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n365_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n407_), .A3(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n413_), .A2(new_n417_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n417_), .B1(new_n413_), .B2(new_n422_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n424_), .A2(new_n425_), .A3(KEYINPUT91), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n413_), .A2(new_n422_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n417_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(KEYINPUT90), .A3(new_n423_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT91), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n362_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n362_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n431_), .B2(KEYINPUT91), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT92), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n437_));
  INV_X1    g236(.A(new_n435_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n426_), .B1(KEYINPUT91), .B2(new_n431_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n437_), .B(new_n438_), .C1(new_n439_), .C2(new_n362_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G22gat), .B(G50gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT93), .ZN(new_n444_));
  INV_X1    g243(.A(G141gat), .ZN(new_n445_));
  INV_X1    g244(.A(G148gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT93), .B1(G141gat), .B2(G148gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(G155gat), .A2(G162gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT1), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G155gat), .A2(G162gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G141gat), .A2(G148gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n449_), .A2(new_n453_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT3), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT2), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n458_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n450_), .A2(new_n452_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n456_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT28), .B1(new_n466_), .B2(KEYINPUT29), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n466_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n443_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n467_), .A3(new_n442_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT96), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G211gat), .B(G218gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(KEYINPUT94), .A2(G197gat), .ZN(new_n479_));
  INV_X1    g278(.A(G204gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(KEYINPUT94), .A2(G197gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT21), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(G197gat), .B2(G204gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n478_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n480_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(G197gat), .A2(G204gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n483_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n479_), .A2(new_n481_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n487_), .B1(new_n490_), .B2(G204gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n477_), .A2(new_n483_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(KEYINPUT95), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT95), .B1(new_n491_), .B2(new_n492_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n489_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n466_), .A2(KEYINPUT29), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G228gat), .A2(G233gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(G78gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(new_n224_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n496_), .A2(new_n497_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n474_), .A2(new_n476_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(new_n476_), .B2(new_n505_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT99), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n466_), .A2(new_n360_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n456_), .B(new_n465_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(KEYINPUT4), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n466_), .A2(new_n360_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n510_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G29gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT100), .B(G85gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT0), .B(G57gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n509_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n523_));
  OR3_X1    g322(.A1(new_n516_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n507_), .A2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G8gat), .B(G36gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G64gat), .B(G92gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n491_), .A2(new_n492_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n535_), .A2(new_n493_), .B1(new_n488_), .B2(new_n485_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n420_), .A2(new_n407_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G226gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT19), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT20), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G169gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n387_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n384_), .B(KEYINPUT97), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n545_), .A2(new_n373_), .B1(new_n394_), .B2(new_n389_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n541_), .B1(new_n496_), .B2(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n537_), .A2(new_n540_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n496_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n541_), .B1(new_n536_), .B2(new_n546_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n540_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n532_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n532_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(new_n540_), .A3(new_n551_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT20), .B1(new_n536_), .B2(new_n546_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n408_), .A2(new_n412_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n536_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n554_), .B(new_n555_), .C1(new_n558_), .C2(new_n540_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(KEYINPUT27), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT102), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n536_), .B1(new_n420_), .B2(new_n407_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT20), .B1(new_n496_), .B2(new_n547_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n562_), .A2(new_n539_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n540_), .B1(new_n537_), .B2(new_n548_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n532_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n559_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT27), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n561_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AOI211_X1 g368(.A(KEYINPUT102), .B(KEYINPUT27), .C1(new_n566_), .C2(new_n559_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n527_), .B(new_n560_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT103), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT101), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT33), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n525_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n513_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n511_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n577_), .A2(new_n521_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n525_), .A2(new_n574_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n566_), .A2(new_n559_), .A3(new_n575_), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n554_), .A2(KEYINPUT32), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n537_), .A2(new_n548_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n539_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n555_), .A3(new_n581_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n583_), .A2(new_n526_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n580_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n573_), .B1(new_n588_), .B2(new_n507_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n476_), .A2(new_n505_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n476_), .A2(new_n505_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(new_n474_), .ZN(new_n592_));
  AOI211_X1 g391(.A(KEYINPUT101), .B(new_n592_), .C1(new_n580_), .C2(new_n587_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n564_), .A2(new_n565_), .A3(new_n532_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n554_), .B1(new_n585_), .B2(new_n555_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n568_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT102), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n567_), .A2(new_n561_), .A3(new_n568_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n527_), .A4(new_n560_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n572_), .A2(new_n594_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n560_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT104), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT104), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n606_), .B(new_n560_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n592_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n526_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n436_), .A2(new_n440_), .A3(new_n609_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n441_), .A2(new_n603_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n338_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n311_), .A2(new_n612_), .A3(new_n312_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n296_), .A2(KEYINPUT81), .A3(new_n338_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT81), .B1(new_n296_), .B2(new_n338_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n613_), .B(new_n614_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n619_), .A2(new_n615_), .B1(new_n612_), .B2(new_n297_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n618_), .B1(new_n620_), .B2(new_n614_), .ZN(new_n621_));
  XOR2_X1   g420(.A(G113gat), .B(G141gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n618_), .B(new_n626_), .C1(new_n620_), .C2(new_n614_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n611_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n354_), .A2(new_n355_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n354_), .A2(new_n631_), .A3(KEYINPUT105), .A4(new_n355_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n609_), .A2(G1gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n588_), .A2(new_n507_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT101), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n588_), .A2(new_n573_), .A3(new_n507_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n642_), .B(new_n643_), .C1(new_n571_), .C2(KEYINPUT103), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n571_), .A2(KEYINPUT103), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n441_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n605_), .A2(new_n607_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n610_), .A3(new_n507_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n280_), .A2(new_n281_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n630_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n330_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n350_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n609_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n640_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n639_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n202_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n662_), .A2(KEYINPUT107), .A3(new_n640_), .A4(new_n658_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(new_n647_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n334_), .B1(new_n656_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n647_), .A2(G8gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n634_), .A2(new_n635_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n634_), .A2(KEYINPUT108), .A3(new_n635_), .A4(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n668_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n668_), .A2(new_n674_), .A3(KEYINPUT40), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n657_), .B2(new_n441_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT41), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n636_), .A2(G15gat), .A3(new_n441_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1326gat));
  OAI21_X1  g482(.A(G22gat), .B1(new_n657_), .B2(new_n507_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT42), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n507_), .A2(G22gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n636_), .B2(new_n686_), .ZN(G1327gat));
  NOR2_X1   g486(.A1(new_n653_), .A2(new_n350_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n652_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G29gat), .B1(new_n689_), .B2(new_n526_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n331_), .A2(new_n352_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n611_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n649_), .A2(new_n694_), .A3(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n350_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n651_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT44), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n701_), .B(new_n698_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n526_), .A2(G29gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n690_), .B1(new_n703_), .B2(new_n704_), .ZN(G1328gat));
  OR2_X1    g504(.A1(new_n665_), .A2(KEYINPUT109), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n665_), .A2(KEYINPUT109), .ZN(new_n707_));
  AOI21_X1  g506(.A(G36gat), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n652_), .A2(new_n708_), .A3(new_n688_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n700_), .A2(new_n702_), .A3(new_n647_), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT46), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n696_), .A2(new_n699_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n701_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n696_), .A2(KEYINPUT44), .A3(new_n699_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n665_), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n711_), .B1(new_n721_), .B2(G36gat), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n722_), .A2(KEYINPUT110), .A3(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n717_), .A2(new_n724_), .ZN(G1329gat));
  INV_X1    g524(.A(new_n441_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n703_), .A2(G43gat), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n689_), .A2(new_n726_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n415_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n689_), .B2(new_n592_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n592_), .A2(G50gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n703_), .B2(new_n734_), .ZN(G1331gat));
  INV_X1    g534(.A(new_n630_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n282_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n649_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(new_n654_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n609_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n738_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n691_), .A2(new_n697_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n609_), .A2(G57gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n706_), .A2(new_n707_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n739_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n747_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n744_), .B2(new_n752_), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n740_), .B2(new_n441_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT49), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n441_), .A2(G71gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n744_), .B2(new_n756_), .ZN(G1334gat));
  OAI21_X1  g556(.A(G78gat), .B1(new_n740_), .B2(new_n507_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT50), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n507_), .A2(G78gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n744_), .B2(new_n760_), .ZN(G1335gat));
  NAND2_X1  g560(.A1(new_n742_), .A2(new_n688_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n211_), .B1(new_n762_), .B2(new_n609_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n764_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n737_), .A2(new_n697_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n696_), .A2(new_n768_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n769_), .A2(new_n211_), .A3(new_n609_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n765_), .A2(new_n766_), .A3(new_n770_), .ZN(G1336gat));
  INV_X1    g570(.A(new_n762_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G92gat), .B1(new_n772_), .B2(new_n665_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n767_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n748_), .A2(new_n210_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT114), .ZN(G1337gat));
  AOI21_X1  g576(.A(new_n234_), .B1(new_n774_), .B2(new_n726_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n726_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n762_), .A2(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n778_), .A2(new_n780_), .A3(KEYINPUT51), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT51), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n778_), .A2(new_n780_), .A3(new_n784_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n787_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n789_), .A2(new_n782_), .A3(KEYINPUT51), .A4(new_n785_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1338gat));
  NAND3_X1  g590(.A1(new_n772_), .A2(new_n224_), .A3(new_n592_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n507_), .B(new_n767_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n224_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n774_), .B2(new_n592_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n793_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n696_), .A2(new_n795_), .A3(new_n592_), .A4(new_n768_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G106gat), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n801_), .A2(KEYINPUT52), .A3(new_n797_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n792_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT53), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n792_), .C1(new_n799_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1339gat));
  OAI21_X1  g606(.A(new_n267_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n264_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n258_), .A2(new_n262_), .A3(new_n267_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT55), .A3(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n274_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n276_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n736_), .A2(new_n277_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n629_), .ZN(new_n822_));
  OAI22_X1  g621(.A1(new_n616_), .A2(new_n617_), .B1(new_n338_), .B2(new_n296_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n626_), .B1(new_n823_), .B2(new_n614_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n614_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n313_), .A2(new_n612_), .B1(new_n619_), .B2(new_n615_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n824_), .A2(new_n825_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n822_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n278_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n330_), .B1(new_n821_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT57), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n811_), .B1(KEYINPUT55), .B2(new_n808_), .ZN(new_n837_));
  AND4_X1   g636(.A1(KEYINPUT55), .A2(new_n259_), .A3(new_n260_), .A4(new_n263_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n816_), .B(new_n274_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n830_), .A2(new_n277_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n816_), .B1(new_n813_), .B2(new_n274_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n843_), .A2(KEYINPUT58), .B1(new_n331_), .B2(new_n352_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n836_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n832_), .A2(new_n835_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n697_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n743_), .A2(new_n851_), .A3(new_n282_), .A4(new_n630_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT54), .B1(new_n353_), .B2(new_n736_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n441_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n608_), .A2(new_n526_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n736_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n855_), .A2(KEYINPUT59), .A3(new_n857_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n736_), .A2(G113gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT121), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n860_), .B1(new_n864_), .B2(new_n866_), .ZN(G1340gat));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n282_), .B2(KEYINPUT60), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n859_), .B(new_n869_), .C1(KEYINPUT60), .C2(new_n868_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n282_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n868_), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n859_), .A2(new_n873_), .A3(new_n350_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n697_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n873_), .ZN(G1342gat));
  AOI21_X1  g675(.A(G134gat), .B1(new_n859_), .B2(new_n330_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT122), .B(G134gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n692_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n864_), .B2(new_n879_), .ZN(G1343gat));
  NAND2_X1  g679(.A1(new_n850_), .A2(new_n854_), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n748_), .A2(new_n726_), .A3(new_n609_), .A4(new_n507_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n630_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n445_), .ZN(G1344gat));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n282_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n446_), .ZN(G1345gat));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n883_), .B2(new_n697_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n881_), .A2(KEYINPUT123), .A3(new_n350_), .A4(new_n882_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n883_), .B2(new_n692_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n653_), .A2(G162gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n883_), .B2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(new_n748_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n898_), .A2(new_n526_), .A3(new_n592_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n832_), .A2(new_n835_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n821_), .A2(new_n831_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n834_), .B1(new_n901_), .B2(new_n330_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n350_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n852_), .A2(new_n853_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n726_), .B(new_n899_), .C1(new_n903_), .C2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT62), .B(G169gat), .C1(new_n905_), .C2(new_n630_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n855_), .A2(new_n736_), .A3(new_n542_), .A4(new_n899_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n881_), .A2(new_n736_), .A3(new_n726_), .A4(new_n899_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT62), .B1(new_n909_), .B2(G169gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT124), .B1(new_n908_), .B2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G169gat), .B1(new_n905_), .B2(new_n630_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n914_), .A2(new_n915_), .A3(new_n906_), .A4(new_n907_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n911_), .A2(new_n916_), .ZN(G1348gat));
  XOR2_X1   g716(.A(KEYINPUT125), .B(G176gat), .Z(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n905_), .A2(new_n282_), .ZN(new_n920_));
  MUX2_X1   g719(.A(new_n918_), .B(new_n919_), .S(new_n920_), .Z(G1349gat));
  NOR2_X1   g720(.A1(new_n905_), .A2(new_n697_), .ZN(new_n922_));
  MUX2_X1   g721(.A(G183gat), .B(new_n390_), .S(new_n922_), .Z(G1350gat));
  OAI21_X1  g722(.A(G190gat), .B1(new_n905_), .B2(new_n692_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n330_), .A2(new_n391_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n905_), .B2(new_n925_), .ZN(G1351gat));
  NAND2_X1  g725(.A1(new_n441_), .A2(new_n527_), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT126), .Z(new_n928_));
  NOR2_X1   g727(.A1(new_n898_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n881_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n736_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n930_), .A2(new_n282_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AND2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  NOR4_X1   g737(.A1(new_n930_), .A2(new_n697_), .A3(new_n937_), .A4(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n931_), .A2(new_n350_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n937_), .ZN(G1354gat));
  OR3_X1    g740(.A1(new_n930_), .A2(G218gat), .A3(new_n653_), .ZN(new_n942_));
  OAI21_X1  g741(.A(G218gat), .B1(new_n930_), .B2(new_n692_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1355gat));
endmodule


