//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n851_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G29gat), .B(G36gat), .Z(new_n210_));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n212_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT76), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G229gat), .A2(G233gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n212_), .B(KEYINPUT15), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n209_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT77), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G169gat), .B(G197gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n228_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n223_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n234_));
  INV_X1    g033(.A(G85gat), .ZN(new_n235_));
  INV_X1    g034(.A(G92gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OR3_X1    g038(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT6), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(G99gat), .B2(G106gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT6), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n240_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT64), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n248_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n239_), .B1(new_n245_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT8), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(KEYINPUT8), .B(new_n239_), .C1(new_n245_), .C2(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n243_), .A2(KEYINPUT6), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n241_), .A2(G99gat), .A3(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n258_));
  INV_X1    g057(.A(G106gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n237_), .A2(KEYINPUT9), .A3(new_n238_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n238_), .A2(KEYINPUT9), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n257_), .A2(new_n261_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G57gat), .B(G64gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G71gat), .B(G78gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT11), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  INV_X1    g067(.A(G64gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G57gat), .ZN(new_n270_));
  INV_X1    g069(.A(G57gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G64gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n272_), .A3(KEYINPUT11), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n265_), .A2(KEYINPUT11), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n267_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n253_), .A2(new_n254_), .A3(new_n264_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G230gat), .A2(G233gat), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n253_), .A2(new_n254_), .A3(new_n264_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n281_));
  INV_X1    g080(.A(new_n276_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n279_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n278_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n277_), .A2(KEYINPUT65), .ZN(new_n288_));
  INV_X1    g087(.A(new_n264_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n254_), .A4(new_n276_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n292_), .A3(KEYINPUT66), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n280_), .A2(new_n282_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT66), .B1(new_n288_), .B2(new_n292_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n287_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(KEYINPUT67), .B(new_n287_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n286_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G120gat), .B(G148gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT69), .ZN(new_n303_));
  XOR2_X1   g102(.A(G176gat), .B(G204gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n234_), .B1(new_n301_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n300_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n288_), .A2(new_n292_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(new_n294_), .A3(new_n293_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT67), .B1(new_n313_), .B2(new_n287_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n285_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n307_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(KEYINPUT70), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n308_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n285_), .B(new_n307_), .C1(new_n309_), .C2(new_n314_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n301_), .A2(KEYINPUT71), .A3(new_n307_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT13), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n323_), .A3(KEYINPUT13), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G226gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT19), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n330_), .B(KEYINPUT89), .Z(new_n331_));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT24), .ZN(new_n333_));
  OR2_X1    g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  MUX2_X1   g133(.A(KEYINPUT24), .B(new_n333_), .S(new_n334_), .Z(new_n335_));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT23), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(G183gat), .A3(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G190gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT25), .B(G183gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT26), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n342_), .B1(new_n345_), .B2(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n335_), .B(new_n340_), .C1(new_n343_), .C2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n337_), .B(KEYINPUT80), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n339_), .B(KEYINPUT81), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT82), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT22), .B(G169gat), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n356_), .A2(KEYINPUT79), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(KEYINPUT79), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n357_), .A2(new_n358_), .B1(G169gat), .B2(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n351_), .A2(KEYINPUT82), .A3(new_n352_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n348_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT85), .B(G197gat), .Z(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(G204gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n366_), .A2(KEYINPUT87), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT21), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n366_), .B2(KEYINPUT87), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT88), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n371_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n366_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n365_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n368_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n364_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(G204gat), .ZN(new_n379_));
  INV_X1    g178(.A(G204gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(G197gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT86), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT21), .B1(new_n379_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n374_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n362_), .A2(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n372_), .A2(new_n373_), .B1(new_n383_), .B2(new_n377_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n351_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n341_), .A2(new_n344_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n335_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n340_), .B1(G183gat), .B2(G190gat), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n356_), .A2(new_n332_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n388_), .A2(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT20), .B1(new_n387_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n331_), .B1(new_n386_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396_));
  INV_X1    g195(.A(new_n393_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n396_), .B1(new_n385_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n362_), .A2(new_n385_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n330_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n387_), .A2(KEYINPUT90), .A3(new_n393_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G64gat), .B(G92gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT92), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n395_), .A2(new_n403_), .A3(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n410_), .A2(KEYINPUT27), .ZN(new_n411_));
  INV_X1    g210(.A(new_n409_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n330_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n400_), .B1(new_n387_), .B2(new_n393_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n399_), .B2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n415_), .A2(KEYINPUT96), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n400_), .B1(new_n385_), .B2(new_n397_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n331_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n417_), .B(new_n418_), .C1(new_n362_), .C2(new_n385_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(new_n415_), .B2(KEYINPUT96), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n412_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n395_), .A2(new_n403_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n412_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n410_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n425_));
  AOI22_X1  g224(.A1(new_n411_), .A2(new_n421_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT2), .ZN(new_n427_));
  INV_X1    g226(.A(G141gat), .ZN(new_n428_));
  INV_X1    g227(.A(G148gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G141gat), .A2(G148gat), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n430_), .B(new_n431_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n435_), .A2(KEYINPUT84), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(KEYINPUT84), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(G155gat), .A2(G162gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G155gat), .A2(G162gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n439_), .B1(KEYINPUT1), .B2(new_n441_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n441_), .A2(KEYINPUT1), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n428_), .A2(new_n429_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n446_), .A2(new_n433_), .A3(new_n447_), .ZN(new_n448_));
  OR3_X1    g247(.A1(new_n443_), .A2(KEYINPUT29), .A3(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n449_), .A2(KEYINPUT28), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(KEYINPUT28), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT29), .B1(new_n443_), .B2(new_n448_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n385_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n385_), .A2(new_n453_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n455_), .A3(new_n451_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G228gat), .A2(G233gat), .ZN(new_n457_));
  INV_X1    g256(.A(G78gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(new_n259_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G22gat), .B(G50gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n454_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n426_), .A2(KEYINPUT99), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n421_), .A2(new_n411_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n410_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n409_), .B1(new_n395_), .B2(new_n403_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n425_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT99), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G225gat), .A2(G233gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(G127gat), .B(G134gat), .Z(new_n476_));
  XOR2_X1   g275(.A(G113gat), .B(G120gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n447_), .A2(new_n433_), .ZN(new_n481_));
  OAI221_X1 g280(.A(new_n478_), .B1(new_n446_), .B2(new_n481_), .C1(new_n438_), .C2(new_n442_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n443_), .A2(new_n448_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(KEYINPUT93), .A3(new_n478_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(KEYINPUT4), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT4), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n480_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n475_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n475_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G1gat), .B(G29gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT94), .B(G85gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT0), .B(G57gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT97), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(KEYINPUT97), .A3(new_n501_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G71gat), .B(G99gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(G43gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(G15gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n507_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n362_), .B(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT83), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n362_), .B(KEYINPUT30), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n511_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n515_), .A2(new_n516_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n511_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n478_), .B(KEYINPUT31), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n518_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n513_), .A2(KEYINPUT83), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n525_), .B2(new_n519_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n514_), .A2(new_n511_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n522_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n504_), .B(new_n505_), .C1(new_n524_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n474_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n524_), .A2(new_n528_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n465_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n467_), .A2(new_n470_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n468_), .A2(new_n469_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT33), .B1(new_n493_), .B2(new_n498_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n493_), .A2(KEYINPUT33), .A3(new_n498_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n491_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n475_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n541_), .A2(new_n498_), .A3(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n537_), .A2(new_n539_), .A3(new_n540_), .A4(new_n543_), .ZN(new_n544_));
  OAI211_X1 g343(.A(KEYINPUT32), .B(new_n409_), .C1(new_n416_), .C2(new_n420_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n395_), .A3(new_n403_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n502_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n533_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n532_), .B1(new_n536_), .B2(new_n551_), .ZN(new_n552_));
  AOI211_X1 g351(.A(new_n233_), .B(new_n328_), .C1(new_n531_), .C2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n221_), .A2(new_n280_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  OAI221_X1 g355(.A(new_n554_), .B1(KEYINPUT35), .B2(new_n556_), .C1(new_n213_), .C2(new_n280_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT72), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n557_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n560_), .A2(KEYINPUT36), .A3(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(KEYINPUT36), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n208_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n282_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT74), .ZN(new_n574_));
  NOR2_X1   g373(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n575_));
  AND2_X1   g374(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n573_), .B(new_n574_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT16), .ZN(new_n579_));
  XOR2_X1   g378(.A(G183gat), .B(G211gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT17), .B1(new_n574_), .B2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n581_), .B1(new_n572_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n573_), .A2(new_n581_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n569_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n553_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n504_), .A2(new_n505_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n203_), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT38), .ZN(new_n592_));
  INV_X1    g391(.A(new_n590_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n328_), .A2(new_n587_), .A3(new_n233_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n567_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n531_), .B2(new_n552_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(KEYINPUT100), .ZN(new_n597_));
  INV_X1    g396(.A(new_n532_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n544_), .A2(new_n550_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n465_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n426_), .A2(new_n504_), .A3(new_n505_), .A4(new_n533_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n598_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n529_), .B1(new_n473_), .B2(new_n466_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n567_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n594_), .B1(new_n597_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n596_), .A2(KEYINPUT100), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n605_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(KEYINPUT101), .A3(new_n594_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n593_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n592_), .B1(new_n203_), .B2(new_n614_), .ZN(G1324gat));
  NAND3_X1  g414(.A1(new_n589_), .A2(new_n204_), .A3(new_n535_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(new_n535_), .A3(new_n594_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n204_), .B1(KEYINPUT102), .B2(KEYINPUT39), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n616_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT40), .B(new_n616_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  NAND3_X1  g425(.A1(new_n589_), .A2(new_n509_), .A3(new_n598_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n612_), .A2(KEYINPUT101), .A3(new_n594_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT101), .B1(new_n612_), .B2(new_n594_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n598_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n630_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT41), .B1(new_n630_), .B2(G15gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n627_), .B1(new_n631_), .B2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n589_), .A2(new_n634_), .A3(new_n533_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n533_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(G22gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n636_), .B2(G22gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(G1327gat));
  INV_X1    g439(.A(new_n587_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(new_n567_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n553_), .A2(new_n642_), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n643_), .A2(G29gat), .A3(new_n593_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n569_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n328_), .A2(new_n233_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT43), .B(new_n569_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n647_), .A2(new_n587_), .A3(new_n648_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n641_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n648_), .A4(new_n649_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n590_), .A3(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n655_), .A2(KEYINPUT103), .A3(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT103), .B1(new_n655_), .B2(G29gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n644_), .B1(new_n656_), .B2(new_n657_), .ZN(G1328gat));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n535_), .A3(new_n654_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G36gat), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n426_), .A2(G36gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n553_), .A2(new_n642_), .A3(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT45), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n660_), .A2(KEYINPUT46), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NAND4_X1  g467(.A1(new_n652_), .A2(G43gat), .A3(new_n598_), .A4(new_n654_), .ZN(new_n669_));
  INV_X1    g468(.A(G43gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n643_), .B2(new_n532_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g472(.A1(new_n652_), .A2(new_n533_), .A3(new_n654_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(G50gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G50gat), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n465_), .A2(G50gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT105), .ZN(new_n679_));
  OAI22_X1  g478(.A1(new_n676_), .A2(new_n677_), .B1(new_n643_), .B2(new_n679_), .ZN(G1331gat));
  AND3_X1   g479(.A1(new_n318_), .A2(new_n323_), .A3(KEYINPUT13), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT13), .B1(new_n318_), .B2(new_n323_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n232_), .B(new_n683_), .C1(new_n531_), .C2(new_n552_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(new_n588_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n271_), .A3(new_n590_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n587_), .A2(new_n232_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n328_), .A2(new_n687_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n612_), .A2(new_n590_), .A3(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n689_), .B2(new_n271_), .ZN(G1332gat));
  NAND3_X1  g489(.A1(new_n685_), .A2(new_n269_), .A3(new_n535_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n612_), .A2(new_n535_), .A3(new_n688_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT48), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G64gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G64gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1333gat));
  INV_X1    g495(.A(G71gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n685_), .A2(new_n697_), .A3(new_n598_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n612_), .A2(new_n598_), .A3(new_n688_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G71gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n702_), .A3(G71gat), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n704_));
  AND3_X1   g503(.A1(new_n701_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n698_), .B1(new_n705_), .B2(new_n706_), .ZN(G1334gat));
  NAND3_X1  g506(.A1(new_n685_), .A2(new_n458_), .A3(new_n533_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n612_), .A2(new_n533_), .A3(new_n688_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT50), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G78gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G78gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1335gat));
  NAND2_X1  g512(.A1(new_n684_), .A2(new_n642_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT108), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n684_), .A2(new_n716_), .A3(new_n642_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n590_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n590_), .A2(G85gat), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT110), .Z(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n683_), .A2(new_n232_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n653_), .A2(new_n649_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n653_), .A2(KEYINPUT109), .A3(new_n649_), .A4(new_n724_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n720_), .A2(KEYINPUT111), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(new_n719_), .B2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1336gat));
  NAND3_X1  g533(.A1(new_n718_), .A2(new_n236_), .A3(new_n535_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n426_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(new_n236_), .ZN(G1337gat));
  AND2_X1   g536(.A1(new_n258_), .A2(new_n260_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n718_), .A2(new_n598_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n532_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n740_));
  INV_X1    g539(.A(G99gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT51), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n739_), .B(new_n744_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1338gat));
  NAND3_X1  g545(.A1(new_n718_), .A2(new_n259_), .A3(new_n533_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n653_), .A2(new_n533_), .A3(new_n649_), .A4(new_n724_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(G106gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G106gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n747_), .B(new_n753_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1339gat));
  AND2_X1   g556(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n758_));
  NOR2_X1   g557(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT113), .B1(new_n683_), .B2(new_n687_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n326_), .A2(KEYINPUT113), .A3(new_n327_), .A4(new_n687_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n567_), .B(new_n568_), .Z(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n761_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n326_), .A2(new_n327_), .A3(new_n687_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n768_), .A2(new_n763_), .A3(new_n758_), .A4(new_n762_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n308_), .A2(new_n317_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n218_), .B1(new_n208_), .B2(new_n212_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n230_), .B1(new_n222_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n217_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n219_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n231_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n771_), .B1(new_n772_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n777_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n324_), .A2(KEYINPUT117), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n319_), .A2(new_n320_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT71), .B1(new_n301_), .B2(new_n307_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT115), .B(new_n232_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n285_), .A2(KEYINPUT55), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n279_), .B(new_n786_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n283_), .A2(new_n284_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n287_), .B1(new_n790_), .B2(new_n310_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n788_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n316_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT56), .B(new_n316_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n784_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT115), .B1(new_n323_), .B2(new_n232_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n567_), .B1(new_n781_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT57), .B(new_n567_), .C1(new_n781_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n798_), .A2(new_n779_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n323_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT118), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n763_), .B1(new_n808_), .B2(KEYINPUT58), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT118), .B(new_n810_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n805_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n770_), .B1(new_n587_), .B2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n474_), .A2(new_n590_), .A3(new_n598_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(G113gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n232_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n815_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n802_), .A2(new_n803_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n641_), .B1(new_n822_), .B2(new_n805_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT59), .B(new_n821_), .C1(new_n823_), .C2(new_n770_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n233_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n818_), .B1(new_n825_), .B2(new_n817_), .ZN(G1340gat));
  AOI21_X1  g625(.A(new_n683_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n827_));
  INV_X1    g626(.A(G120gat), .ZN(new_n828_));
  INV_X1    g627(.A(new_n816_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(KEYINPUT60), .B2(new_n828_), .ZN(new_n831_));
  OAI22_X1  g630(.A1(new_n827_), .A2(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n816_), .B2(new_n641_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n820_), .A2(new_n824_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n641_), .A2(G127gat), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT119), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n833_), .B1(new_n834_), .B2(new_n836_), .ZN(G1342gat));
  INV_X1    g636(.A(G134gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n816_), .A2(new_n838_), .A3(new_n595_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n763_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n838_), .ZN(G1343gat));
  NOR4_X1   g640(.A1(new_n593_), .A2(new_n598_), .A3(new_n535_), .A4(new_n465_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT120), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n813_), .A2(new_n587_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n770_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n232_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n328_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT121), .B(G148gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1345gat));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n641_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1346gat));
  INV_X1    g654(.A(G162gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n847_), .B2(new_n569_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n595_), .A2(new_n856_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n814_), .A2(new_n844_), .A3(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT122), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n847_), .A2(new_n856_), .A3(new_n595_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n569_), .B(new_n843_), .C1(new_n823_), .C2(new_n770_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G162gat), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n865_), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n529_), .A2(new_n426_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n232_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT123), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n465_), .B(new_n869_), .C1(new_n823_), .C2(new_n770_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n870_), .A2(G169gat), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n870_), .B2(G169gat), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n465_), .B(new_n867_), .C1(new_n823_), .C2(new_n770_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n232_), .A2(new_n354_), .ZN(new_n875_));
  OAI22_X1  g674(.A1(new_n872_), .A2(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1348gat));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n683_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(G176gat), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n874_), .A2(new_n355_), .A3(new_n683_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1349gat));
  NOR2_X1   g679(.A1(new_n874_), .A2(new_n587_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(G183gat), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n874_), .A2(new_n344_), .A3(new_n587_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n874_), .B2(new_n763_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n595_), .A2(new_n341_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n874_), .B2(new_n886_), .ZN(G1351gat));
  NAND3_X1  g686(.A1(new_n532_), .A2(new_n593_), .A3(new_n533_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n889_), .A2(KEYINPUT125), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(KEYINPUT125), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n535_), .A3(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n814_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(G197gat), .A4(new_n232_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n892_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n232_), .B(new_n896_), .C1(new_n823_), .C2(new_n770_), .ZN(new_n897_));
  INV_X1    g696(.A(G197gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT126), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n898_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n895_), .A2(new_n899_), .A3(new_n900_), .ZN(G1352gat));
  NAND2_X1  g700(.A1(new_n893_), .A2(new_n328_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G204gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n893_), .A2(new_n380_), .A3(new_n328_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1353gat));
  OAI211_X1 g704(.A(new_n641_), .B(new_n896_), .C1(new_n823_), .C2(new_n770_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AND2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n906_), .B2(new_n907_), .ZN(G1354gat));
  NAND2_X1  g709(.A1(new_n893_), .A2(new_n595_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT127), .B(G218gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n763_), .A2(new_n912_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n911_), .A2(new_n912_), .B1(new_n893_), .B2(new_n913_), .ZN(G1355gat));
endmodule


