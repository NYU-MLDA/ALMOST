//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G71gat), .B(G78gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n205_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n207_), .B1(new_n210_), .B2(new_n206_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT64), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT65), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n215_), .A2(new_n217_), .A3(new_n222_), .A4(new_n218_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n220_), .A2(KEYINPUT67), .A3(new_n221_), .A4(new_n223_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT6), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n212_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n212_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .A4(new_n229_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n232_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT8), .B1(new_n233_), .B2(KEYINPUT66), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n231_), .A2(KEYINPUT8), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT10), .B(G99gat), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n214_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT9), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(G85gat), .A3(G92gat), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n239_), .A2(new_n241_), .A3(new_n229_), .A4(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n211_), .B1(new_n238_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n211_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n234_), .A2(new_n235_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n248_), .A2(new_n212_), .A3(new_n237_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT8), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n224_), .A2(new_n225_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n229_), .A3(new_n227_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n252_), .B2(new_n212_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n244_), .B(new_n247_), .C1(new_n249_), .C2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n246_), .A2(KEYINPUT12), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n256_), .B(new_n211_), .C1(new_n238_), .C2(new_n245_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n203_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  AOI211_X1 g057(.A(KEYINPUT68), .B(new_n202_), .C1(new_n246_), .C2(new_n254_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n246_), .A2(new_n254_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT68), .B1(new_n261_), .B2(new_n202_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT5), .B(G176gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G120gat), .B(G148gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n260_), .A2(new_n262_), .A3(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n268_), .A2(KEYINPUT13), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT13), .B1(new_n268_), .B2(new_n270_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G29gat), .B(G36gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G43gat), .B(G50gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n276_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n274_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G15gat), .B(G22gat), .ZN(new_n283_));
  INV_X1    g082(.A(G1gat), .ZN(new_n284_));
  INV_X1    g083(.A(G8gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT14), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G8gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n287_), .B(new_n288_), .Z(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT74), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n282_), .A2(new_n289_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G229gat), .A3(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n280_), .B(KEYINPUT15), .ZN(new_n295_));
  INV_X1    g094(.A(new_n289_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G229gat), .A2(G233gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n290_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G113gat), .B(G141gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G169gat), .B(G197gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n303_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n294_), .A2(new_n299_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n273_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT104), .ZN(new_n311_));
  XOR2_X1   g110(.A(G141gat), .B(G148gat), .Z(new_n312_));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT81), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(G155gat), .A3(G162gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n312_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OR3_X1    g122(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n324_), .A2(new_n326_), .A3(new_n327_), .A4(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n314_), .A2(new_n316_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(new_n320_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n323_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(KEYINPUT29), .ZN(new_n333_));
  XOR2_X1   g132(.A(G22gat), .B(G50gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(G204gat), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT21), .ZN(new_n341_));
  INV_X1    g140(.A(G197gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(G204gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT87), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G211gat), .B(G218gat), .Z(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n342_), .ZN(new_n350_));
  INV_X1    g149(.A(G204gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n342_), .A2(G204gat), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n350_), .A2(KEYINPUT86), .A3(new_n351_), .A4(new_n352_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n348_), .B1(new_n358_), .B2(KEYINPUT21), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n340_), .A2(new_n344_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n341_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n348_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n340_), .A2(new_n344_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(KEYINPUT88), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n347_), .A2(new_n359_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT83), .B(G228gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT84), .B(G233gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n366_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n370_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n358_), .A2(KEYINPUT21), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n345_), .A2(KEYINPUT87), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n360_), .A2(new_n346_), .A3(new_n341_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n376_), .A2(new_n363_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n362_), .A2(new_n365_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT89), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n379_), .A2(new_n380_), .B1(new_n372_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n322_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(new_n320_), .A3(new_n318_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n328_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n327_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(new_n325_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n319_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n384_), .A2(new_n312_), .B1(new_n390_), .B2(new_n330_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT89), .B1(new_n391_), .B2(new_n371_), .ZN(new_n392_));
  AOI211_X1 g191(.A(KEYINPUT90), .B(new_n375_), .C1(new_n382_), .C2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n379_), .A2(new_n380_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n372_), .A2(new_n381_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n392_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n397_), .B2(new_n370_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n374_), .B1(new_n393_), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n381_), .B1(new_n332_), .B2(KEYINPUT29), .ZN(new_n403_));
  AOI211_X1 g202(.A(KEYINPUT89), .B(new_n371_), .C1(new_n323_), .C2(new_n331_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n366_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT90), .B1(new_n405_), .B2(new_n375_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n394_), .A3(new_n370_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(new_n374_), .A3(new_n400_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n402_), .A2(KEYINPUT91), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT91), .B1(new_n402_), .B2(new_n409_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n337_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT19), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT94), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G183gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT25), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT76), .B(G190gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT26), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G169gat), .ZN(new_n428_));
  INV_X1    g227(.A(G176gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(KEYINPUT24), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G183gat), .A2(G190gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT23), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n425_), .B(KEYINPUT77), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT24), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n424_), .A2(new_n432_), .A3(new_n434_), .A4(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(G176gat), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OR3_X1    g240(.A1(new_n441_), .A2(KEYINPUT78), .A3(new_n430_), .ZN(new_n442_));
  INV_X1    g241(.A(G183gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n421_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n434_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT78), .B1(new_n441_), .B2(new_n430_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n438_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n415_), .B1(new_n366_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n438_), .A2(new_n447_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n395_), .A2(KEYINPUT94), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT22), .B(G169gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n439_), .A2(KEYINPUT92), .A3(new_n440_), .ZN(new_n456_));
  AOI21_X1  g255(.A(G176gat), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT93), .B1(new_n457_), .B2(new_n430_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n456_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT92), .B1(new_n439_), .B2(new_n440_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n429_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT93), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n431_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n434_), .B1(G183gat), .B2(G190gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT26), .B(G190gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT25), .B(G183gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n432_), .A2(new_n437_), .A3(new_n434_), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT20), .B1(new_n470_), .B2(new_n395_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n414_), .B1(new_n452_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n395_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n414_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n366_), .A2(new_n448_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n473_), .A2(KEYINPUT20), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478_));
  INV_X1    g277(.A(G92gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT18), .B(G64gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n465_), .A2(new_n469_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n366_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n487_), .A2(new_n474_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n473_), .A2(KEYINPUT20), .A3(new_n475_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n414_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n490_), .A3(new_n482_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n484_), .A2(KEYINPUT27), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT27), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n488_), .A2(new_n490_), .A3(new_n482_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n482_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n400_), .B1(new_n408_), .B2(new_n374_), .ZN(new_n499_));
  AOI211_X1 g298(.A(new_n373_), .B(new_n401_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n337_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n412_), .A2(new_n497_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT80), .B(G127gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(G113gat), .A2(G120gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G113gat), .A2(G120gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(G134gat), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(G134gat), .B1(new_n507_), .B2(new_n508_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n506_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n511_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n509_), .A3(new_n505_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n323_), .A2(new_n512_), .A3(new_n514_), .A4(new_n331_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n323_), .A2(new_n331_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n512_), .A2(new_n514_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n332_), .A2(KEYINPUT95), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT4), .B1(new_n519_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT96), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G225gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n332_), .A2(new_n520_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n527_), .A2(KEYINPUT4), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT97), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n516_), .A3(new_n515_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n521_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT96), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT4), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .A4(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT98), .B1(new_n531_), .B2(new_n525_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n537_));
  XNOR2_X1  g336(.A(G1gat), .B(G29gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G85gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n532_), .B1(new_n531_), .B2(KEYINPUT4), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544_));
  AOI211_X1 g343(.A(KEYINPUT96), .B(new_n544_), .C1(new_n530_), .C2(new_n521_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n546_), .A2(KEYINPUT98), .A3(new_n526_), .A4(new_n529_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n536_), .A2(new_n542_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n542_), .B1(new_n536_), .B2(new_n547_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G227gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n520_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(new_n448_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n448_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G71gat), .B(G99gat), .ZN(new_n557_));
  INV_X1    g356(.A(G43gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(KEYINPUT30), .B(G15gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n555_), .A2(new_n556_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n550_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n311_), .B1(new_n504_), .B2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n402_), .A2(new_n409_), .A3(KEYINPUT91), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n502_), .B1(new_n501_), .B2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n411_), .A2(new_n337_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n564_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n571_), .A2(KEYINPUT104), .A3(new_n572_), .A4(new_n497_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n567_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n549_), .A2(KEYINPUT33), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT33), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n576_), .B(new_n542_), .C1(new_n536_), .C2(new_n547_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n495_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n546_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n541_), .B1(new_n531_), .B2(new_n526_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT100), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n578_), .B(new_n491_), .C1(new_n579_), .C2(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n575_), .A2(new_n577_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT102), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n482_), .A2(KEYINPUT32), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n477_), .B2(new_n586_), .ZN(new_n587_));
  AOI211_X1 g386(.A(KEYINPUT102), .B(new_n585_), .C1(new_n472_), .C2(new_n476_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n585_), .B(KEYINPUT101), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n488_), .A2(new_n490_), .A3(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n589_), .B(new_n591_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n571_), .B1(new_n583_), .B2(new_n593_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n550_), .B(new_n497_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT103), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n412_), .A2(new_n503_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n598_), .A2(KEYINPUT103), .A3(new_n550_), .A4(new_n497_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n594_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n574_), .B1(new_n600_), .B2(new_n564_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n310_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G162gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT71), .B(G134gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n238_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n244_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n295_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT70), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(KEYINPUT35), .A3(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(KEYINPUT35), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT69), .ZN(new_n617_));
  INV_X1    g416(.A(new_n280_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n610_), .B2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n609_), .A2(KEYINPUT69), .A3(new_n280_), .A4(new_n244_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n611_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n615_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT35), .ZN(new_n624_));
  INV_X1    g423(.A(new_n614_), .ZN(new_n625_));
  AOI211_X1 g424(.A(new_n624_), .B(new_n625_), .C1(new_n611_), .C2(KEYINPUT70), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT36), .B(new_n608_), .C1(new_n622_), .C2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n622_), .A2(new_n627_), .A3(new_n630_), .A4(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n603_), .B1(new_n628_), .B2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(new_n627_), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n629_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(KEYINPUT37), .A3(new_n632_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n289_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(new_n247_), .ZN(new_n641_));
  XOR2_X1   g440(.A(G127gat), .B(G155gat), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(G211gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT16), .B(G183gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n643_), .B(new_n644_), .Z(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT17), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT72), .Z(new_n648_));
  NOR2_X1   g447(.A1(new_n641_), .A2(new_n646_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(KEYINPUT17), .B2(new_n645_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n638_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n602_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT105), .ZN(new_n654_));
  INV_X1    g453(.A(new_n550_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n284_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT38), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n636_), .A2(KEYINPUT106), .A3(new_n632_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT106), .B1(new_n636_), .B2(new_n632_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n651_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n602_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n550_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n657_), .A2(new_n664_), .ZN(G1324gat));
  INV_X1    g464(.A(new_n497_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n654_), .A2(new_n285_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G8gat), .B1(new_n663_), .B2(new_n497_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(KEYINPUT39), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(KEYINPUT39), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(G1325gat));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n662_), .B2(new_n565_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT41), .ZN(new_n676_));
  INV_X1    g475(.A(new_n653_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n674_), .A3(new_n565_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1326gat));
  INV_X1    g478(.A(G22gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n662_), .B2(new_n598_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT42), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n677_), .A2(new_n680_), .A3(new_n598_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1327gat));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n597_), .A2(new_n599_), .ZN(new_n686_));
  OR3_X1    g485(.A1(new_n575_), .A2(new_n577_), .A3(new_n582_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n598_), .B1(new_n687_), .B2(new_n592_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n564_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n574_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n691_), .B2(new_n638_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n638_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n601_), .A2(KEYINPUT43), .A3(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n309_), .B(new_n651_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n691_), .A2(new_n685_), .A3(new_n638_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n601_), .B2(new_n693_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n310_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n651_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702_), .B2(new_n550_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n658_), .A2(new_n659_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n651_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n602_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n550_), .A2(G29gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT107), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n703_), .A2(new_n710_), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n697_), .A2(new_n666_), .A3(new_n701_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n697_), .A2(new_n701_), .A3(KEYINPUT108), .A4(new_n666_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(G36gat), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(KEYINPUT46), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n497_), .B(KEYINPUT109), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n707_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT45), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n716_), .A2(new_n718_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n718_), .B1(new_n716_), .B2(new_n722_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  OAI21_X1  g524(.A(G43gat), .B1(new_n702_), .B2(new_n564_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n707_), .A2(new_n558_), .A3(new_n565_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(G1330gat));
  OAI21_X1  g529(.A(G50gat), .B1(new_n702_), .B2(new_n571_), .ZN(new_n731_));
  INV_X1    g530(.A(G50gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n707_), .A2(new_n732_), .A3(new_n598_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1331gat));
  NOR2_X1   g533(.A1(new_n271_), .A2(new_n272_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(new_n307_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n601_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(new_n652_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G57gat), .B1(new_n739_), .B2(new_n655_), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT111), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n661_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n655_), .B2(KEYINPUT111), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n740_), .B1(new_n742_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(new_n720_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G64gat), .B1(new_n743_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT48), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(G64gat), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT112), .Z(new_n751_));
  NAND2_X1  g550(.A1(new_n739_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n743_), .B2(new_n564_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT49), .ZN(new_n755_));
  INV_X1    g554(.A(G71gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n739_), .A2(new_n756_), .A3(new_n565_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1334gat));
  OAI21_X1  g557(.A(G78gat), .B1(new_n743_), .B2(new_n571_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT50), .ZN(new_n760_));
  INV_X1    g559(.A(G78gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n739_), .A2(new_n761_), .A3(new_n598_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1335gat));
  AND2_X1   g562(.A1(new_n738_), .A2(new_n706_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764_), .B2(new_n655_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n737_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n651_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n550_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n765_), .B1(new_n768_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g568(.A(G92gat), .B1(new_n764_), .B2(new_n666_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n767_), .A2(new_n479_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n720_), .ZN(G1337gat));
  NAND3_X1  g571(.A1(new_n766_), .A2(new_n565_), .A3(new_n651_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n565_), .A2(new_n240_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n773_), .A2(G99gat), .B1(new_n764_), .B2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n777_), .B(new_n778_), .Z(G1338gat));
  NAND3_X1  g578(.A1(new_n764_), .A2(new_n214_), .A3(new_n598_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n766_), .A2(new_n598_), .A3(new_n651_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g585(.A1(new_n634_), .A2(new_n308_), .A3(new_n705_), .A4(new_n637_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n788_), .A2(new_n735_), .A3(new_n790_), .A4(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n791_), .B(new_n792_), .C1(new_n787_), .C2(new_n273_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n255_), .A2(new_n257_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n202_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n259_), .ZN(new_n800_));
  AND4_X1   g599(.A1(new_n262_), .A2(new_n799_), .A3(new_n800_), .A4(new_n269_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n308_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n799_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n255_), .A2(new_n203_), .A3(new_n257_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n258_), .A2(KEYINPUT55), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n267_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT115), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n812_), .B(KEYINPUT56), .C1(new_n808_), .C2(new_n267_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT55), .B1(new_n798_), .B2(new_n202_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n804_), .B(new_n203_), .C1(new_n255_), .C2(new_n257_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n269_), .B1(new_n818_), .B2(new_n806_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n815_), .B1(new_n819_), .B2(KEYINPUT56), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n808_), .A2(new_n815_), .A3(KEYINPUT56), .A4(new_n267_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n803_), .B1(new_n814_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n293_), .A2(new_n298_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n290_), .A2(new_n297_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n825_), .B(new_n303_), .C1(new_n298_), .C2(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n827_), .A2(new_n306_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n269_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n801_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT117), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(new_n828_), .C1(new_n801_), .C2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT57), .B(new_n704_), .C1(new_n824_), .C2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n812_), .B1(new_n819_), .B2(KEYINPUT56), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n267_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT116), .ZN(new_n839_));
  INV_X1    g638(.A(new_n806_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n816_), .A2(new_n817_), .A3(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT115), .B(new_n810_), .C1(new_n841_), .C2(new_n269_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n837_), .A2(new_n839_), .A3(new_n821_), .A4(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n834_), .B1(new_n843_), .B2(new_n802_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n836_), .B1(new_n844_), .B2(new_n660_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n809_), .A2(new_n810_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n838_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n270_), .A3(new_n828_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n847_), .A2(KEYINPUT58), .A3(new_n270_), .A4(new_n828_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n638_), .A3(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n835_), .A2(new_n845_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n797_), .B1(new_n853_), .B2(new_n651_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n550_), .A2(new_n564_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n854_), .A2(new_n504_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G113gat), .B1(new_n857_), .B2(new_n307_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n651_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n797_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n504_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n855_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n866_));
  NAND4_X1  g665(.A1(new_n861_), .A2(new_n862_), .A3(new_n855_), .A4(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n308_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n858_), .B1(new_n868_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g668(.A(G120gat), .ZN(new_n870_));
  INV_X1    g669(.A(new_n864_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n857_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n872_), .B2(new_n273_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n870_), .A2(KEYINPUT60), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n875_));
  AOI21_X1  g674(.A(G120gat), .B1(new_n273_), .B2(new_n875_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n863_), .A2(new_n874_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT119), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879_));
  INV_X1    g678(.A(new_n877_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n735_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n879_), .B(new_n880_), .C1(new_n881_), .C2(new_n870_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n882_), .ZN(G1341gat));
  AOI21_X1  g682(.A(G127gat), .B1(new_n857_), .B2(new_n705_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n651_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g685(.A(G134gat), .B1(new_n857_), .B2(new_n660_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n693_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(G134gat), .ZN(G1343gat));
  NOR4_X1   g688(.A1(new_n720_), .A2(new_n550_), .A3(new_n565_), .A4(new_n571_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT120), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n861_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n308_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT121), .B(G141gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  INV_X1    g694(.A(new_n892_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n273_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g697(.A1(new_n892_), .A2(G155gat), .A3(new_n651_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G155gat), .B1(new_n892_), .B2(new_n651_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n896_), .B2(new_n660_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n638_), .A2(G162gat), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT123), .Z(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n896_), .B2(new_n906_), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n854_), .A2(new_n747_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n598_), .A2(new_n566_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT62), .B(G169gat), .C1(new_n910_), .C2(new_n308_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  INV_X1    g711(.A(new_n909_), .ZN(new_n913_));
  NOR4_X1   g712(.A1(new_n854_), .A2(new_n308_), .A3(new_n747_), .A4(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n914_), .B2(new_n428_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n460_), .B2(new_n459_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT124), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n911_), .A2(new_n915_), .A3(new_n916_), .A4(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1348gat));
  NOR2_X1   g720(.A1(new_n910_), .A2(new_n735_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n429_), .ZN(G1349gat));
  NOR2_X1   g722(.A1(new_n910_), .A2(new_n651_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n467_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n443_), .B2(new_n924_), .ZN(G1350gat));
  NAND4_X1  g725(.A1(new_n908_), .A2(new_n466_), .A3(new_n660_), .A4(new_n909_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n861_), .A2(new_n638_), .A3(new_n720_), .A4(new_n909_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n928_), .A2(new_n929_), .A3(G190gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n928_), .B2(G190gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n927_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT126), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n934_), .B(new_n927_), .C1(new_n930_), .C2(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1351gat));
  NAND2_X1  g735(.A1(new_n598_), .A2(new_n550_), .ZN(new_n937_));
  NOR4_X1   g736(.A1(new_n854_), .A2(new_n565_), .A3(new_n937_), .A4(new_n747_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n307_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n273_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n705_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n943_), .B2(new_n944_), .ZN(G1354gat));
  INV_X1    g746(.A(G218gat), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n938_), .A2(new_n948_), .A3(new_n660_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n948_), .B1(new_n938_), .B2(new_n638_), .ZN(new_n951_));
  OAI21_X1  g750(.A(KEYINPUT127), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n938_), .A2(new_n638_), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n953_), .B(new_n949_), .C1(new_n954_), .C2(new_n948_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n952_), .A2(new_n955_), .ZN(G1355gat));
endmodule


