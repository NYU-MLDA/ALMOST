//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G218gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G211gat), .ZN(new_n206_));
  INV_X1    g005(.A(G211gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G218gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT87), .ZN(new_n211_));
  INV_X1    g010(.A(G204gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(G197gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT21), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(KEYINPUT87), .B2(new_n202_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(G197gat), .ZN(new_n216_));
  INV_X1    g015(.A(G197gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G204gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n206_), .B(new_n208_), .C1(new_n219_), .C2(KEYINPUT21), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n210_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n221_), .A2(KEYINPUT86), .B1(G228gat), .B2(G233gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n209_), .B1(new_n203_), .B2(new_n202_), .ZN(new_n224_));
  OAI211_X1 g023(.A(KEYINPUT21), .B(new_n213_), .C1(new_n219_), .C2(new_n211_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n224_), .A2(new_n225_), .B1(new_n209_), .B2(new_n204_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228_));
  INV_X1    g027(.A(G141gat), .ZN(new_n229_));
  INV_X1    g028(.A(G148gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT2), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n231_), .A2(new_n234_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n243_), .A3(new_n239_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n239_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT1), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n229_), .A2(new_n230_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n244_), .A2(new_n246_), .A3(new_n232_), .A4(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n227_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(G78gat), .B1(new_n226_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(new_n248_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT29), .ZN(new_n252_));
  INV_X1    g051(.A(G78gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n221_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n254_), .A3(G106gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(G106gat), .B1(new_n250_), .B2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n223_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G22gat), .B(G50gat), .Z(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n251_), .B2(KEYINPUT29), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n251_), .A2(KEYINPUT29), .A3(new_n261_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n260_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G106gat), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n226_), .A2(new_n249_), .A3(G78gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n253_), .B1(new_n252_), .B2(new_n221_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(new_n222_), .A3(new_n255_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n258_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n267_), .A3(KEYINPUT88), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT89), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT89), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n265_), .A2(new_n267_), .A3(KEYINPUT88), .A4(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n276_), .A2(new_n281_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT90), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT80), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n292_), .A4(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G183gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT25), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G183gat), .ZN(new_n298_));
  INV_X1    g097(.A(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT26), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G190gat), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n296_), .A2(new_n298_), .A3(new_n300_), .A4(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n294_), .A2(new_n303_), .A3(new_n307_), .A4(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT83), .B(G176gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT22), .B(G169gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n306_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n295_), .A2(new_n299_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n304_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n316_), .A3(new_n292_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n310_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n287_), .B1(new_n318_), .B2(new_n226_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n316_), .A2(new_n292_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT22), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n289_), .A2(KEYINPUT81), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT81), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G169gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT82), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT82), .B1(new_n321_), .B2(G169gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n311_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n320_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n291_), .A2(new_n293_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n308_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n333_), .A2(new_n294_), .A3(new_n307_), .A4(new_n303_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n334_), .A3(new_n226_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n310_), .A2(new_n317_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n221_), .A2(new_n336_), .A3(KEYINPUT90), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n319_), .A2(KEYINPUT20), .A3(new_n335_), .A4(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT19), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n226_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT20), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n221_), .B2(new_n336_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n342_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n345_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n318_), .B2(new_n226_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n316_), .A2(new_n292_), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT83), .B(G176gat), .Z(new_n351_));
  NOR2_X1   g150(.A1(new_n323_), .A2(G169gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n289_), .A2(KEYINPUT81), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT22), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n329_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n351_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n350_), .B1(new_n356_), .B2(new_n327_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n334_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n221_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n349_), .A2(new_n359_), .A3(KEYINPUT91), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n347_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G8gat), .B(G36gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n341_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n341_), .B2(new_n361_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n286_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT20), .B1(new_n221_), .B2(new_n336_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n340_), .B1(new_n343_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n365_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n341_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT27), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n368_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n285_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n331_), .A2(new_n334_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT30), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT84), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381_));
  INV_X1    g180(.A(G43gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384_));
  INV_X1    g183(.A(G15gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n383_), .B(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n380_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n379_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G134gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G127gat), .ZN(new_n393_));
  INV_X1    g192(.A(G127gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G134gat), .ZN(new_n395_));
  INV_X1    g194(.A(G120gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G113gat), .ZN(new_n397_));
  INV_X1    g196(.A(G113gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G120gat), .ZN(new_n399_));
  AND4_X1   g198(.A1(new_n393_), .A2(new_n395_), .A3(new_n397_), .A4(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n393_), .A2(new_n395_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT31), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OR3_X1    g203(.A1(new_n388_), .A2(new_n391_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(G85gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT0), .B(G57gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n251_), .A2(new_n412_), .A3(new_n402_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n417_));
  INV_X1    g216(.A(new_n236_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n235_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n240_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n245_), .A2(new_n425_), .A3(KEYINPUT1), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n247_), .B(new_n232_), .C1(new_n243_), .C2(new_n239_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n402_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n242_), .B(new_n248_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(KEYINPUT92), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT92), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n251_), .A2(new_n432_), .A3(new_n402_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n417_), .B1(new_n434_), .B2(KEYINPUT4), .ZN(new_n435_));
  AOI211_X1 g234(.A(KEYINPUT93), .B(new_n412_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n416_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n414_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n411_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT97), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AOI211_X1 g240(.A(KEYINPUT97), .B(new_n411_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n438_), .A2(new_n411_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n441_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n377_), .A2(new_n407_), .A3(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n368_), .B(new_n375_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT33), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n366_), .A2(new_n367_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n413_), .A2(new_n414_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n411_), .B1(new_n434_), .B2(new_n415_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n452_), .A2(new_n453_), .A3(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n438_), .A2(KEYINPUT33), .A3(new_n411_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n437_), .A2(KEYINPUT94), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT94), .B1(new_n437_), .B2(new_n459_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT95), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT96), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n341_), .A2(new_n361_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n464_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n341_), .A2(new_n361_), .A3(KEYINPUT96), .A4(new_n466_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n468_), .A2(new_n469_), .B1(new_n467_), .B2(new_n371_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n445_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n470_), .B1(new_n471_), .B2(new_n442_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n437_), .A2(new_n459_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n437_), .A2(KEYINPUT94), .A3(new_n459_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n465_), .A2(new_n372_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n457_), .A2(new_n374_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n477_), .A2(new_n479_), .A3(new_n480_), .A4(new_n452_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n463_), .A2(new_n472_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n450_), .B1(new_n482_), .B2(new_n284_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n448_), .B1(new_n483_), .B2(new_n407_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT73), .B(G1gat), .ZN(new_n485_));
  INV_X1    g284(.A(G8gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G8gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G29gat), .B(G36gat), .Z(new_n495_));
  XOR2_X1   g294(.A(G43gat), .B(G50gat), .Z(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  XOR2_X1   g296(.A(new_n494_), .B(new_n497_), .Z(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G229gat), .A3(G233gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n494_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(new_n497_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT78), .Z(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G169gat), .B(G197gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT79), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n508_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n484_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n517_));
  OR2_X1    g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n521_));
  OR2_X1    g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT10), .B(G99gat), .Z(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(G99gat), .A3(G106gat), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n524_), .A2(new_n271_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n522_), .A2(new_n523_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT66), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n271_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT7), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n528_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n531_), .A2(new_n536_), .A3(new_n532_), .A4(new_n271_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT8), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT67), .ZN(new_n540_));
  INV_X1    g339(.A(new_n519_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n518_), .A2(KEYINPUT67), .A3(new_n519_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n538_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n539_), .B1(new_n538_), .B2(new_n545_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n530_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G57gat), .B(G64gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT11), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G78gat), .Z(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n549_), .A2(KEYINPUT11), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(KEYINPUT12), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT69), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT69), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n548_), .A2(new_n558_), .A3(KEYINPUT12), .A4(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT64), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT12), .B1(new_n548_), .B2(new_n555_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n548_), .A2(new_n555_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT68), .B1(new_n548_), .B2(new_n555_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n555_), .B2(new_n548_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT68), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n569_), .B(new_n562_), .C1(new_n570_), .C2(new_n565_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n567_), .A2(new_n571_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(KEYINPUT13), .A3(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT70), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n582_), .A2(KEYINPUT70), .A3(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n548_), .A2(new_n497_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT72), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n501_), .A2(new_n548_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n592_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(KEYINPUT36), .ZN(new_n603_));
  INV_X1    g402(.A(new_n598_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n591_), .A2(new_n604_), .A3(new_n596_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n599_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n602_), .B(KEYINPUT36), .Z(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n599_), .B2(new_n605_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n606_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n599_), .A2(new_n605_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n607_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n599_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n610_), .A2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n555_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n494_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(KEYINPUT76), .ZN(new_n620_));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT75), .ZN(new_n622_));
  XOR2_X1   g421(.A(G127gat), .B(G155gat), .Z(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n618_), .B(new_n502_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT17), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n626_), .A2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n620_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n619_), .A2(KEYINPUT76), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n628_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n619_), .A2(KEYINPUT17), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n632_), .B(new_n633_), .C1(new_n634_), .C2(new_n626_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n631_), .A2(new_n635_), .A3(KEYINPUT77), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT77), .B1(new_n631_), .B2(new_n635_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n616_), .A2(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n516_), .A2(new_n589_), .A3(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n446_), .A3(new_n485_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT38), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT99), .B1(new_n606_), .B2(new_n609_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n612_), .A2(new_n645_), .A3(new_n614_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n484_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n631_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n635_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n588_), .A2(new_n514_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n648_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n447_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n641_), .A2(new_n642_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n643_), .A2(new_n655_), .A3(new_n656_), .ZN(G1324gat));
  NAND3_X1  g456(.A1(new_n648_), .A2(new_n376_), .A3(new_n653_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G8gat), .B1(new_n658_), .B2(new_n659_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n661_), .A2(new_n662_), .A3(KEYINPUT39), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT39), .B1(new_n661_), .B2(new_n662_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n640_), .A2(new_n486_), .A3(new_n376_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(KEYINPUT40), .A3(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  INV_X1    g470(.A(new_n407_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G15gat), .B1(new_n654_), .B2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT41), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n640_), .A2(new_n385_), .A3(new_n407_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n654_), .B2(new_n284_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n640_), .A2(new_n679_), .A3(new_n285_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1327gat));
  INV_X1    g480(.A(new_n638_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n588_), .A2(new_n682_), .A3(new_n647_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n516_), .A2(new_n683_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n684_), .A2(G29gat), .A3(new_n447_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n638_), .A2(new_n586_), .A3(new_n515_), .A4(new_n587_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT101), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n484_), .A2(new_n688_), .A3(new_n616_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n484_), .B2(new_n616_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n687_), .B(KEYINPUT44), .C1(new_n689_), .C2(new_n690_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n446_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(new_n696_), .A3(G29gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(G29gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n685_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT103), .B(new_n685_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n693_), .A2(new_n376_), .A3(new_n694_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n376_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n516_), .A2(new_n683_), .A3(new_n708_), .ZN(new_n709_));
  XOR2_X1   g508(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n704_), .B1(new_n706_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1329gat));
  NOR2_X1   g513(.A1(new_n672_), .A2(new_n382_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n693_), .A2(new_n694_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT106), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n693_), .A2(new_n718_), .A3(new_n694_), .A4(new_n715_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n382_), .B1(new_n684_), .B2(new_n672_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(G1330gat));
  OR3_X1    g522(.A1(new_n684_), .A2(G50gat), .A3(new_n284_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n693_), .A2(KEYINPUT108), .A3(new_n285_), .A4(new_n694_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(G50gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n693_), .A2(new_n285_), .A3(new_n694_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n725_), .B1(new_n727_), .B2(new_n730_), .ZN(new_n731_));
  AND4_X1   g530(.A1(new_n725_), .A2(new_n730_), .A3(G50gat), .A4(new_n726_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n724_), .B1(new_n731_), .B2(new_n732_), .ZN(G1331gat));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n484_), .A2(new_n734_), .A3(new_n514_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n484_), .B2(new_n514_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n639_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n737_), .A2(new_n589_), .A3(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n446_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n514_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n589_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n648_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n447_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n741_), .A2(new_n746_), .ZN(G1332gat));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n744_), .B2(new_n376_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT48), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n748_), .A3(new_n376_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n744_), .B2(new_n407_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT49), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n739_), .A2(new_n753_), .A3(new_n407_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1334gat));
  AOI21_X1  g556(.A(new_n253_), .B1(new_n744_), .B2(new_n285_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT50), .Z(new_n759_));
  NAND3_X1  g558(.A1(new_n739_), .A2(new_n253_), .A3(new_n285_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1335gat));
  NOR3_X1   g560(.A1(new_n589_), .A2(new_n682_), .A3(new_n647_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT111), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n762_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G85gat), .B1(new_n767_), .B2(new_n446_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n689_), .A2(new_n690_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n589_), .A2(new_n515_), .A3(new_n682_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n446_), .A2(G85gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT112), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n768_), .B1(new_n772_), .B2(new_n774_), .ZN(G1336gat));
  INV_X1    g574(.A(G92gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n767_), .A2(new_n776_), .A3(new_n376_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n772_), .A2(new_n376_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n779_), .B2(new_n776_), .ZN(G1337gat));
  NAND3_X1  g579(.A1(new_n767_), .A2(new_n407_), .A3(new_n524_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G99gat), .B1(new_n771_), .B2(new_n672_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n781_), .B(new_n782_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n784_), .B2(KEYINPUT113), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(G1338gat));
  OAI211_X1 g586(.A(new_n285_), .B(new_n770_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G106gat), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT52), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n284_), .A2(G106gat), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n767_), .A2(KEYINPUT115), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT115), .B1(new_n767_), .B2(new_n791_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n790_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n616_), .A2(new_n742_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n584_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NOR4_X1   g601(.A1(new_n616_), .A2(new_n742_), .A3(new_n584_), .A4(KEYINPUT54), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n610_), .A2(new_n615_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n579_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n512_), .B1(new_n499_), .B2(new_n507_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n498_), .A2(new_n506_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n506_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n503_), .A2(new_n504_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n511_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n807_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n806_), .A2(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n560_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT116), .B1(new_n814_), .B2(KEYINPUT55), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n563_), .B1(new_n560_), .B2(new_n566_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n814_), .B2(KEYINPUT55), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n567_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n576_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n576_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n813_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n805_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT58), .B(new_n813_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n514_), .A2(new_n806_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n812_), .B1(new_n579_), .B2(new_n577_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n829_), .B1(new_n834_), .B2(new_n647_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n644_), .A2(new_n646_), .ZN(new_n836_));
  AOI211_X1 g635(.A(KEYINPUT57), .B(new_n836_), .C1(new_n831_), .C2(new_n833_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n828_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n804_), .B1(new_n838_), .B2(new_n652_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n377_), .A2(new_n407_), .A3(new_n446_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n804_), .B1(new_n838_), .B2(new_n638_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n844_), .A2(KEYINPUT59), .A3(new_n840_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n398_), .A2(KEYINPUT117), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n398_), .B1(new_n515_), .B2(KEYINPUT117), .ZN(new_n847_));
  NOR4_X1   g646(.A1(new_n843_), .A2(new_n845_), .A3(new_n846_), .A4(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G113gat), .B1(new_n841_), .B2(new_n515_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT118), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n843_), .A2(new_n845_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n847_), .A2(new_n846_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854_));
  INV_X1    g653(.A(new_n849_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n850_), .A2(new_n856_), .ZN(G1340gat));
  INV_X1    g656(.A(new_n851_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G120gat), .B1(new_n858_), .B2(new_n589_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860_));
  AOI21_X1  g659(.A(G120gat), .B1(new_n588_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT119), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n860_), .B2(G120gat), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n841_), .B(new_n862_), .C1(new_n861_), .C2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n859_), .A2(new_n865_), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n858_), .B2(new_n652_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n841_), .A2(new_n394_), .A3(new_n682_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1342gat));
  OAI21_X1  g668(.A(G134gat), .B1(new_n858_), .B2(new_n805_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n841_), .A2(new_n392_), .A3(new_n836_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1343gat));
  NAND4_X1  g671(.A1(new_n672_), .A2(new_n285_), .A3(new_n446_), .A4(new_n707_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n839_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n515_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n588_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT120), .B(G148gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1345gat));
  NAND2_X1  g678(.A1(new_n874_), .A2(new_n682_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  AOI21_X1  g681(.A(G162gat), .B1(new_n874_), .B2(new_n836_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT121), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n616_), .A2(G162gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n874_), .B2(new_n885_), .ZN(G1347gat));
  NOR3_X1   g685(.A1(new_n672_), .A2(new_n446_), .A3(new_n707_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n284_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n844_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n289_), .B1(new_n889_), .B2(new_n515_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n890_), .A2(KEYINPUT62), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n312_), .A3(new_n515_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(KEYINPUT62), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(G1348gat));
  AOI21_X1  g693(.A(new_n351_), .B1(new_n889_), .B2(new_n588_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n839_), .A2(new_n285_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n887_), .A2(new_n588_), .A3(G176gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1349gat));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n682_), .A3(new_n887_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n652_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n899_), .A2(new_n295_), .B1(new_n889_), .B2(new_n900_), .ZN(G1350gat));
  NAND4_X1  g700(.A1(new_n889_), .A2(new_n300_), .A3(new_n302_), .A4(new_n836_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n844_), .A2(new_n805_), .A3(new_n888_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n299_), .ZN(G1351gat));
  NOR4_X1   g703(.A1(new_n407_), .A2(new_n446_), .A3(new_n284_), .A4(new_n707_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n839_), .A2(KEYINPUT122), .A3(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n800_), .A2(new_n801_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT54), .ZN(new_n910_));
  INV_X1    g709(.A(new_n803_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n830_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n914_));
  INV_X1    g713(.A(new_n820_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n560_), .A2(KEYINPUT55), .A3(new_n563_), .A4(new_n566_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n557_), .A2(new_n559_), .B1(new_n565_), .B2(new_n564_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n563_), .B2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n818_), .B1(new_n567_), .B2(new_n819_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n915_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n914_), .B1(new_n920_), .B2(new_n578_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n576_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n913_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n647_), .B1(new_n923_), .B2(new_n832_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT57), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n834_), .A2(new_n829_), .A3(new_n647_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n925_), .A2(new_n926_), .B1(new_n827_), .B2(new_n826_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n912_), .B1(new_n927_), .B2(new_n651_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n908_), .B1(new_n928_), .B2(new_n905_), .ZN(new_n929_));
  OAI211_X1 g728(.A(G197gat), .B(new_n515_), .C1(new_n907_), .C2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT122), .B1(new_n839_), .B2(new_n906_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n928_), .A2(new_n908_), .A3(new_n905_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n935_), .A2(KEYINPUT123), .A3(G197gat), .A4(new_n515_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n932_), .A2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n515_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n217_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT124), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n938_), .A2(new_n941_), .A3(new_n217_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n937_), .B1(new_n940_), .B2(new_n942_), .ZN(G1352gat));
  INV_X1    g742(.A(new_n935_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n589_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(new_n212_), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT125), .B(G204gat), .Z(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n945_), .B2(new_n948_), .ZN(G1353gat));
  AOI211_X1 g748(.A(KEYINPUT63), .B(G211gat), .C1(new_n935_), .C2(new_n651_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n944_), .A2(new_n652_), .ZN(new_n951_));
  XOR2_X1   g750(.A(KEYINPUT63), .B(G211gat), .Z(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(G1354gat));
  AOI21_X1  g752(.A(G218gat), .B1(new_n935_), .B2(new_n836_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n805_), .A2(new_n205_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(KEYINPUT126), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n935_), .B2(new_n956_), .ZN(G1355gat));
endmodule


