//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT65), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT9), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n208_), .A2(new_n209_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n212_), .B(new_n213_), .C1(new_n211_), .C2(KEYINPUT9), .ZN(new_n214_));
  INV_X1    g013(.A(new_n213_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n215_), .A2(new_n211_), .A3(KEYINPUT9), .A4(new_n210_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n205_), .A2(new_n207_), .A3(new_n214_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT67), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n207_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n215_), .A2(new_n210_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(KEYINPUT8), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(KEYINPUT8), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n217_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G78gat), .Z(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n217_), .B(new_n234_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G230gat), .A2(G233gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT64), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n242_), .A2(KEYINPUT68), .ZN(new_n243_));
  INV_X1    g042(.A(new_n237_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(new_n236_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n227_), .A2(KEYINPUT12), .A3(new_n235_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n247_), .A2(KEYINPUT69), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(KEYINPUT69), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n240_), .B(new_n246_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(KEYINPUT68), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n243_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G120gat), .B(G148gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G176gat), .B(G204gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n243_), .A2(new_n250_), .A3(new_n251_), .A4(new_n258_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT13), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT13), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n252_), .A2(new_n258_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n260_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G231gat), .A2(G233gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n234_), .B(new_n268_), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT73), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271_));
  INV_X1    g070(.A(G1gat), .ZN(new_n272_));
  INV_X1    g071(.A(G8gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT14), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G1gat), .B(G8gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n270_), .B(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G127gat), .B(G155gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(G183gat), .B(G211gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT17), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n278_), .A2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n284_), .A2(KEYINPUT17), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n278_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G29gat), .B(G36gat), .Z(new_n290_));
  XOR2_X1   g089(.A(G43gat), .B(G50gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT15), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n227_), .A2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n295_));
  NAND2_X1  g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT35), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT72), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n292_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n294_), .B(new_n299_), .C1(new_n300_), .C2(new_n227_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n297_), .A2(new_n298_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G190gat), .B(G218gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G134gat), .B(G162gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT36), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n308_), .B(KEYINPUT36), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT37), .B1(new_n311_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n305_), .A2(new_n312_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT37), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n316_), .B(new_n317_), .C1(new_n310_), .C2(new_n305_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n289_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n267_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT75), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n293_), .A2(new_n277_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n300_), .A2(new_n277_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G229gat), .A2(G233gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n300_), .B(new_n277_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G113gat), .B(G141gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT76), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G169gat), .B(G197gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  OR2_X1    g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n325_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338_));
  INV_X1    g137(.A(G169gat), .ZN(new_n339_));
  INV_X1    g138(.A(G176gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT78), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348_));
  INV_X1    g147(.A(G183gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(KEYINPUT77), .A2(G183gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT25), .A3(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n349_), .A2(KEYINPUT25), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT26), .B(G190gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n341_), .A2(new_n344_), .A3(new_n356_), .A4(new_n345_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n347_), .A2(new_n355_), .A3(new_n357_), .A4(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362_));
  NOR2_X1   g161(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G169gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n350_), .A2(new_n351_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(G190gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n344_), .A2(new_n345_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n361_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n362_), .B1(new_n361_), .B2(new_n368_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G15gat), .B(G43gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT81), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n373_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(G71gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G99gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n374_), .A2(new_n375_), .A3(new_n383_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(KEYINPUT83), .A3(new_n386_), .ZN(new_n390_));
  INV_X1    g189(.A(G134gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G127gat), .ZN(new_n392_));
  INV_X1    g191(.A(G127gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(G134gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G120gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G113gat), .ZN(new_n397_));
  INV_X1    g196(.A(G113gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G120gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n392_), .A2(new_n394_), .A3(new_n397_), .A4(new_n399_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n395_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n405_), .A2(KEYINPUT82), .A3(new_n397_), .A4(new_n399_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT31), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n389_), .A2(new_n390_), .A3(new_n408_), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n387_), .A2(new_n388_), .A3(new_n408_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G197gat), .B(G204gat), .Z(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT21), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G211gat), .B(G218gat), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G197gat), .B(G204gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT21), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(new_n418_), .A3(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G155gat), .B(G162gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G141gat), .A2(G148gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT2), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n422_), .A2(KEYINPUT85), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n422_), .B2(KEYINPUT85), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT84), .B1(new_n429_), .B2(KEYINPUT3), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G141gat), .A2(G148gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT3), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n421_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n421_), .A2(KEYINPUT1), .ZN(new_n437_));
  NAND3_X1  g236(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n429_), .A2(new_n422_), .A3(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT29), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n420_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G22gat), .B(G50gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n442_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT87), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G228gat), .A2(G233gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n450_), .B(G78gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(new_n204_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(new_n448_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n449_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n445_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n457_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n445_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n455_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n407_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n421_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n425_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n422_), .A2(KEYINPUT85), .A3(new_n423_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n426_), .ZN(new_n467_));
  NOR4_X1   g266(.A1(KEYINPUT84), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n432_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n464_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n440_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n401_), .A2(new_n403_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G225gat), .A2(G233gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n463_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n463_), .A2(KEYINPUT4), .A3(new_n474_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n475_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n463_), .B2(KEYINPUT4), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT89), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n471_), .A2(new_n472_), .B1(new_n406_), .B2(new_n404_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT4), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n475_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n463_), .A2(KEYINPUT4), .A3(new_n474_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n481_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n476_), .B1(new_n480_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G1gat), .B(G29gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(G85gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT0), .B(G57gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT89), .B1(new_n477_), .B2(new_n479_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n484_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n476_), .A2(new_n491_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT93), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n500_));
  AOI211_X1 g299(.A(new_n500_), .B(new_n497_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n493_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G8gat), .B(G36gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT18), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G64gat), .B(G92gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT32), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G226gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT19), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT20), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n349_), .A2(KEYINPUT25), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n354_), .A2(new_n353_), .A3(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n344_), .A2(new_n345_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n514_), .A2(new_n360_), .A3(new_n515_), .A4(new_n341_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(G183gat), .A2(G190gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n364_), .B1(new_n367_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n512_), .B1(new_n420_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n361_), .A2(new_n368_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT79), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n361_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n511_), .B(new_n520_), .C1(new_n524_), .C2(new_n420_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n420_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n415_), .A2(new_n419_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n519_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n512_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n511_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n525_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AOI211_X1 g331(.A(KEYINPUT91), .B(new_n511_), .C1(new_n526_), .C2(new_n529_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n508_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT92), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n369_), .A2(new_n370_), .A3(new_n420_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n520_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n510_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n526_), .A2(new_n511_), .A3(new_n529_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n536_), .B1(new_n541_), .B2(new_n508_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n539_), .A2(KEYINPUT90), .A3(new_n540_), .A4(new_n507_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT20), .B1(new_n420_), .B2(new_n519_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n524_), .B2(new_n420_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT91), .B1(new_n546_), .B2(new_n511_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n530_), .A2(new_n531_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n525_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n508_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n502_), .A2(new_n535_), .A3(new_n544_), .A4(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n498_), .B1(new_n480_), .B2(new_n486_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT33), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT33), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n496_), .A2(new_n555_), .A3(new_n498_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n539_), .A2(new_n506_), .A3(new_n540_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n506_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT88), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n485_), .B(new_n475_), .C1(KEYINPUT4), .C2(new_n463_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n463_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n492_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n506_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n541_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n558_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n557_), .A2(new_n561_), .A3(new_n564_), .A4(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n462_), .B1(new_n552_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n506_), .B(KEYINPUT94), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n549_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(KEYINPUT27), .A3(new_n558_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT27), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n553_), .A2(new_n500_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n496_), .A2(KEYINPUT93), .A3(new_n498_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n462_), .A2(new_n579_), .A3(new_n493_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n411_), .B1(new_n570_), .B2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n409_), .A2(new_n410_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n502_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n462_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n576_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .A4(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n337_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n321_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n584_), .A2(G1gat), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT38), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT96), .Z(new_n592_));
  NOR3_X1   g391(.A1(new_n266_), .A2(new_n337_), .A3(new_n289_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n311_), .A2(new_n314_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n272_), .B1(new_n597_), .B2(new_n502_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n589_), .A2(KEYINPUT38), .A3(new_n590_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT95), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(KEYINPUT95), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n598_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n592_), .A2(new_n602_), .ZN(G1324gat));
  NAND3_X1  g402(.A1(new_n589_), .A2(new_n273_), .A3(new_n576_), .ZN(new_n604_));
  AOI211_X1 g403(.A(KEYINPUT39), .B(new_n273_), .C1(new_n597_), .C2(new_n576_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n597_), .A2(new_n576_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n607_), .B2(G8gat), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n596_), .B2(new_n411_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT41), .Z(new_n612_));
  INV_X1    g411(.A(new_n589_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n411_), .A2(G15gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(G1326gat));
  OAI21_X1  g414(.A(G22gat), .B1(new_n596_), .B2(new_n585_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT42), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n585_), .A2(G22gat), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n613_), .B2(new_n618_), .ZN(G1327gat));
  INV_X1    g418(.A(new_n594_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n289_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n266_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(new_n588_), .ZN(new_n623_));
  AOI21_X1  g422(.A(G29gat), .B1(new_n623_), .B2(new_n502_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n266_), .A2(new_n337_), .A3(new_n621_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT43), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n582_), .A2(new_n587_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n315_), .A2(new_n318_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n626_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT43), .B(new_n628_), .C1(new_n582_), .C2(new_n587_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n625_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  OAI211_X1 g434(.A(KEYINPUT97), .B(new_n625_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n267_), .A2(new_n336_), .A3(new_n289_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n627_), .A2(new_n629_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT43), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n627_), .A2(new_n626_), .A3(new_n629_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT44), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n637_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n502_), .A2(G29gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n624_), .B1(new_n645_), .B2(new_n646_), .ZN(G1328gat));
  INV_X1    g446(.A(G36gat), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n576_), .A2(KEYINPUT99), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n576_), .A2(KEYINPUT99), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n623_), .A2(new_n648_), .A3(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(KEYINPUT100), .B(KEYINPUT45), .Z(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT101), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n652_), .B(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n586_), .B1(new_n642_), .B2(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n637_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n658_), .B2(G36gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT98), .B(new_n648_), .C1(new_n637_), .C2(new_n657_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT46), .B(new_n655_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1329gat));
  INV_X1    g464(.A(G43gat), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n411_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT102), .B1(new_n644_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n637_), .A2(new_n643_), .A3(new_n670_), .A4(new_n667_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n623_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n672_), .B2(new_n411_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT47), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n669_), .A2(new_n676_), .A3(new_n671_), .A4(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n623_), .B2(new_n462_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n462_), .A2(G50gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n645_), .B2(new_n680_), .ZN(G1331gat));
  NAND2_X1  g480(.A1(new_n266_), .A2(new_n337_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n319_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT103), .Z(new_n685_));
  NOR2_X1   g484(.A1(new_n584_), .A2(G57gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n682_), .A2(new_n289_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n595_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n502_), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n685_), .A2(new_n686_), .B1(G57gat), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(G1332gat));
  INV_X1    g492(.A(new_n651_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G64gat), .B1(new_n688_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT48), .ZN(new_n696_));
  INV_X1    g495(.A(new_n685_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n694_), .A2(G64gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n697_), .B2(new_n698_), .ZN(G1333gat));
  NOR3_X1   g498(.A1(new_n697_), .A2(G71gat), .A3(new_n411_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n689_), .A2(new_n583_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G71gat), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT105), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n701_), .A2(new_n704_), .A3(G71gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT49), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n703_), .A2(KEYINPUT49), .A3(new_n705_), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n700_), .A2(new_n706_), .A3(new_n707_), .ZN(G1334gat));
  OAI21_X1  g507(.A(G78gat), .B1(new_n688_), .B2(new_n585_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT50), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n585_), .A2(G78gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n697_), .B2(new_n711_), .ZN(G1335gat));
  NAND2_X1  g511(.A1(new_n640_), .A2(new_n641_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n682_), .A2(new_n621_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G85gat), .B1(new_n715_), .B2(new_n584_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n621_), .A2(new_n620_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n683_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n502_), .A2(new_n208_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n716_), .B1(new_n718_), .B2(new_n719_), .ZN(G1336gat));
  OAI21_X1  g519(.A(G92gat), .B1(new_n715_), .B2(new_n694_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n576_), .A2(new_n209_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n718_), .B2(new_n722_), .ZN(G1337gat));
  NAND4_X1  g522(.A1(new_n683_), .A2(new_n583_), .A3(new_n203_), .A4(new_n717_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT106), .ZN(new_n725_));
  OAI21_X1  g524(.A(G99gat), .B1(new_n715_), .B2(new_n411_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(KEYINPUT108), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n727_), .A2(new_n729_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT107), .B1(new_n725_), .B2(new_n726_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(G1338gat));
  XNOR2_X1  g532(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n734_));
  OAI21_X1  g533(.A(G106gat), .B1(new_n715_), .B2(new_n585_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT110), .B(G106gat), .C1(new_n715_), .C2(new_n585_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n736_), .A3(new_n734_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n683_), .A2(new_n204_), .A3(new_n462_), .A4(new_n717_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n739_), .A2(new_n744_), .A3(new_n740_), .A4(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1339gat));
  INV_X1    g545(.A(KEYINPUT57), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n250_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n246_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n241_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n247_), .B(KEYINPUT69), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n752_), .A2(KEYINPUT55), .A3(new_n240_), .A4(new_n246_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n257_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(KEYINPUT56), .A3(new_n257_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n260_), .A2(new_n336_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n260_), .A2(KEYINPUT111), .A3(new_n336_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n259_), .A2(new_n260_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n322_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n333_), .B1(new_n326_), .B2(new_n324_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n335_), .A2(new_n767_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT112), .Z(new_n769_));
  AOI22_X1  g568(.A1(new_n758_), .A2(new_n763_), .B1(new_n764_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n747_), .B1(new_n770_), .B2(new_n594_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n757_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n761_), .B(new_n762_), .C1(new_n772_), .C2(new_n755_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n764_), .A2(new_n769_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT57), .A3(new_n620_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n260_), .B(new_n769_), .C1(new_n772_), .C2(new_n755_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n758_), .A2(KEYINPUT58), .A3(new_n260_), .A4(new_n769_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n629_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n771_), .A2(new_n776_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n289_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n319_), .A2(new_n337_), .A3(new_n265_), .A4(new_n261_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  NOR4_X1   g587(.A1(new_n411_), .A2(new_n576_), .A3(new_n584_), .A4(new_n462_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT116), .B(G113gat), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n337_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n776_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n771_), .A2(new_n781_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(KEYINPUT115), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n771_), .A2(new_n797_), .A3(new_n781_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n621_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n786_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT114), .B(KEYINPUT59), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n789_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n791_), .B(new_n793_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n398_), .B1(new_n790_), .B2(new_n337_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT113), .B(new_n398_), .C1(new_n790_), .C2(new_n337_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n803_), .A2(new_n806_), .A3(new_n807_), .ZN(G1340gat));
  OAI211_X1 g607(.A(new_n266_), .B(new_n791_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n809_));
  XOR2_X1   g608(.A(KEYINPUT117), .B(G120gat), .Z(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n267_), .B2(KEYINPUT60), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(KEYINPUT60), .B2(new_n810_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n790_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(G1341gat));
  NOR2_X1   g615(.A1(new_n289_), .A2(new_n393_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n791_), .B(new_n817_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n393_), .B1(new_n790_), .B2(new_n289_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT118), .B(new_n393_), .C1(new_n790_), .C2(new_n289_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n818_), .A2(new_n821_), .A3(new_n822_), .ZN(G1342gat));
  OAI211_X1 g622(.A(new_n629_), .B(new_n791_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G134gat), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n788_), .A2(new_n391_), .A3(new_n594_), .A4(new_n789_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1343gat));
  AOI21_X1  g626(.A(new_n786_), .B1(new_n782_), .B2(new_n289_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n651_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n828_), .A2(new_n583_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n336_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n266_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g634(.A(KEYINPUT61), .B(G155gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n831_), .A2(new_n838_), .A3(new_n621_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n831_), .B2(new_n621_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n837_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n828_), .A2(new_n583_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n829_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT119), .B1(new_n844_), .B2(new_n289_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n839_), .A3(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(G1346gat));
  INV_X1    g646(.A(G162gat), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n844_), .A2(new_n848_), .A3(new_n628_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n844_), .B2(new_n620_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT120), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n852_), .B(new_n848_), .C1(new_n844_), .C2(new_n620_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n851_), .B2(new_n853_), .ZN(G1347gat));
  NAND3_X1  g653(.A1(new_n651_), .A2(new_n584_), .A3(new_n583_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n462_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n336_), .B(new_n856_), .C1(new_n799_), .C2(new_n786_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT22), .B(G169gat), .Z(new_n858_));
  OR2_X1    g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(KEYINPUT122), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n339_), .B1(new_n860_), .B2(KEYINPUT122), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n857_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n857_), .B2(new_n862_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n859_), .B1(new_n863_), .B2(new_n864_), .ZN(G1348gat));
  OR2_X1    g664(.A1(new_n799_), .A2(new_n786_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n266_), .A3(new_n856_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n828_), .A2(new_n462_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n267_), .A2(new_n855_), .A3(new_n340_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n867_), .A2(new_n340_), .B1(new_n868_), .B2(new_n869_), .ZN(G1349gat));
  NOR2_X1   g669(.A1(new_n855_), .A2(new_n289_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n365_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n289_), .B1(new_n353_), .B2(new_n513_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n856_), .B(new_n873_), .C1(new_n799_), .C2(new_n786_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n872_), .B1(new_n875_), .B2(new_n876_), .ZN(G1350gat));
  NAND3_X1  g676(.A1(new_n866_), .A2(new_n629_), .A3(new_n856_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G190gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n594_), .A2(new_n354_), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT124), .Z(new_n881_));
  NAND3_X1  g680(.A1(new_n866_), .A2(new_n856_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1351gat));
  NOR2_X1   g682(.A1(new_n694_), .A2(new_n580_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n843_), .A2(new_n336_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT126), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n887_), .B(new_n889_), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n843_), .A2(new_n884_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n267_), .ZN(new_n892_));
  AND2_X1   g691(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n892_), .B2(new_n894_), .ZN(G1353gat));
  NAND3_X1  g695(.A1(new_n843_), .A2(new_n621_), .A3(new_n884_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  AND2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n897_), .B2(new_n898_), .ZN(G1354gat));
  OAI21_X1  g700(.A(G218gat), .B1(new_n891_), .B2(new_n628_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n620_), .A2(G218gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n891_), .B2(new_n903_), .ZN(G1355gat));
endmodule


