//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(KEYINPUT77), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT24), .B1(new_n205_), .B2(new_n206_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n210_), .B(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n213_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n205_), .A2(KEYINPUT24), .A3(new_n206_), .A4(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n220_), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT25), .B1(new_n220_), .B2(KEYINPUT75), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n212_), .A2(new_n217_), .A3(new_n219_), .A4(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n211_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n228_));
  OR3_X1    g027(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G227gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(G71gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G99gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT80), .B1(new_n242_), .B2(KEYINPUT79), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n244_), .B(new_n245_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n240_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G113gat), .B(G120gat), .Z(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n243_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n239_), .A2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n237_), .B(new_n238_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G15gat), .B(G43gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT78), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT30), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT31), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n253_), .A2(new_n259_), .A3(new_n254_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT84), .ZN(new_n264_));
  OR2_X1    g063(.A1(G197gat), .A2(G204gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G197gat), .A2(G204gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(KEYINPUT83), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G211gat), .B(G218gat), .Z(new_n272_));
  OAI21_X1  g071(.A(new_n269_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n264_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n271_), .A2(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n272_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(KEYINPUT84), .A3(new_n277_), .A4(new_n269_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n225_), .A2(new_n230_), .A3(new_n275_), .A4(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT20), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT22), .B(G169gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n204_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n218_), .B(KEYINPUT85), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n227_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT25), .B(G183gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n222_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n209_), .A2(new_n211_), .A3(new_n286_), .A4(new_n219_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n273_), .A2(new_n274_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n280_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n279_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT19), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n275_), .A2(new_n278_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n231_), .A2(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n284_), .A2(new_n287_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n289_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n280_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n293_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G8gat), .B(G36gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT18), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n294_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT90), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n294_), .A2(new_n301_), .A3(KEYINPUT90), .A4(new_n305_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n225_), .A2(new_n230_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT20), .B1(new_n288_), .B2(new_n289_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n293_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n279_), .A2(new_n290_), .A3(new_n300_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n305_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(new_n309_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT27), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n310_), .A2(new_n311_), .A3(new_n293_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n300_), .B1(new_n279_), .B2(new_n290_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n315_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT27), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n306_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(KEYINPUT1), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(KEYINPUT81), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n326_), .A2(KEYINPUT1), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n328_), .B2(KEYINPUT81), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT2), .B1(new_n334_), .B2(KEYINPUT82), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n333_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n338_), .A2(new_n341_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n327_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(new_n326_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n337_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n345_), .A2(new_n347_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n336_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT86), .B1(new_n249_), .B2(new_n242_), .ZN(new_n355_));
  OR3_X1    g154(.A1(new_n249_), .A2(KEYINPUT86), .A3(new_n242_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n350_), .A2(new_n357_), .A3(KEYINPUT4), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT87), .B(KEYINPUT4), .Z(new_n361_));
  OAI211_X1 g160(.A(new_n349_), .B(new_n361_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n350_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G85gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT0), .B(G57gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n363_), .A2(new_n364_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT28), .B1(new_n349_), .B2(KEYINPUT29), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT28), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n354_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n376_), .B1(new_n337_), .B2(new_n348_), .ZN(new_n384_));
  OAI211_X1 g183(.A(G228gat), .B(G233gat), .C1(new_n384_), .C2(new_n298_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n295_), .B(new_n386_), .C1(new_n354_), .C2(new_n376_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G22gat), .B(G50gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n383_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n385_), .A2(new_n387_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n388_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n395_), .A2(new_n382_), .A3(new_n380_), .A4(new_n390_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n373_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n325_), .A2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n393_), .A2(new_n396_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n372_), .A2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n321_), .A2(new_n306_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n350_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT88), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n369_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n405_), .B2(new_n369_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n404_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n363_), .A2(KEYINPUT33), .A3(new_n364_), .A4(new_n371_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n402_), .A2(new_n403_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n305_), .A2(KEYINPUT32), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n319_), .A2(new_n320_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n412_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n372_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n371_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n400_), .B1(new_n411_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n399_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI211_X1 g220(.A(KEYINPUT89), .B(new_n400_), .C1(new_n418_), .C2(new_n411_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n263_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n400_), .B1(new_n318_), .B2(new_n324_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n261_), .A2(new_n370_), .A3(new_n262_), .A4(new_n372_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT91), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n429_), .A3(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n423_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT71), .B(G1gat), .ZN(new_n433_));
  INV_X1    g232(.A(G8gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G15gat), .B(G22gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G8gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G29gat), .B(G36gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT67), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n442_), .A2(KEYINPUT67), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n444_), .A2(KEYINPUT68), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT68), .ZN(new_n447_));
  XOR2_X1   g246(.A(G29gat), .B(G36gat), .Z(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n447_), .B1(new_n450_), .B2(new_n443_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G43gat), .B(G50gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n446_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT68), .B1(new_n444_), .B2(new_n445_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n447_), .A3(new_n443_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n441_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n453_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT15), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n440_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n460_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(new_n439_), .ZN(new_n466_));
  OR3_X1    g265(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n465_), .B(new_n439_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n464_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G113gat), .B(G141gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G169gat), .B(G197gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n470_), .B(new_n471_), .Z(new_n472_));
  NAND3_X1  g271(.A1(new_n467_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT66), .B(KEYINPUT34), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G232gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT35), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n458_), .A2(new_n461_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT10), .B(G99gat), .Z(new_n491_));
  INV_X1    g290(.A(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT64), .ZN(new_n495_));
  INV_X1    g294(.A(G85gat), .ZN(new_n496_));
  INV_X1    g295(.A(G92gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT9), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n490_), .B(new_n493_), .C1(new_n495_), .C2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n235_), .A2(new_n492_), .A3(KEYINPUT65), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT7), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n506_), .A2(new_n235_), .A3(new_n492_), .A4(KEYINPUT65), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n490_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT8), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n498_), .A2(new_n500_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n503_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n485_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n481_), .A2(new_n482_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n465_), .B2(new_n513_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n484_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n513_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n520_), .A2(new_n516_), .A3(new_n483_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n478_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G190gat), .B(G218gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT69), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G134gat), .B(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT36), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n528_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n527_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n522_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  OAI221_X1 g331(.A(new_n478_), .B1(new_n532_), .B2(new_n528_), .C1(new_n518_), .C2(new_n521_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n531_), .A2(KEYINPUT37), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT37), .B1(new_n531_), .B2(new_n533_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G127gat), .B(G155gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G183gat), .B(G211gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n542_), .A2(KEYINPUT73), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n546_));
  XOR2_X1   g345(.A(G71gat), .B(G78gat), .Z(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n547_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n552_), .B(KEYINPUT72), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n551_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n439_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI211_X1 g355(.A(new_n544_), .B(new_n556_), .C1(new_n542_), .C2(new_n541_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n555_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n536_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n551_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n513_), .A2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n551_), .B(new_n503_), .C1(new_n512_), .C2(new_n511_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n562_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(KEYINPUT12), .A3(new_n565_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n513_), .A2(new_n568_), .A3(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n566_), .B1(new_n570_), .B2(new_n562_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n576_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n577_), .A2(KEYINPUT13), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT13), .B1(new_n577_), .B2(new_n578_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n432_), .A2(new_n477_), .A3(new_n561_), .A4(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT92), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n433_), .A3(new_n373_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n531_), .A2(new_n533_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT94), .ZN(new_n587_));
  INV_X1    g386(.A(new_n581_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(new_n476_), .ZN(new_n589_));
  AND4_X1   g388(.A1(new_n432_), .A2(new_n559_), .A3(new_n587_), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n373_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n584_), .A2(new_n585_), .B1(G1gat), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n584_), .A2(new_n585_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT93), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT93), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n592_), .B1(new_n594_), .B2(new_n595_), .ZN(G1324gat));
  AOI21_X1  g395(.A(new_n323_), .B1(new_n317_), .B2(KEYINPUT27), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n583_), .A2(new_n434_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n590_), .A2(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(G8gat), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n600_), .A2(KEYINPUT39), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(KEYINPUT39), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n598_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g403(.A(G15gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n263_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n590_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT41), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n583_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1326gat));
  INV_X1    g409(.A(G22gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n590_), .B2(new_n400_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT42), .Z(new_n613_));
  NAND3_X1  g412(.A1(new_n583_), .A2(new_n611_), .A3(new_n400_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1327gat));
  AOI21_X1  g414(.A(new_n429_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n616_));
  NOR4_X1   g415(.A1(new_n597_), .A2(new_n425_), .A3(new_n400_), .A4(KEYINPUT91), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n411_), .A2(new_n418_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT89), .B1(new_n619_), .B2(new_n400_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n419_), .A2(new_n420_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(new_n399_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n618_), .B1(new_n622_), .B2(new_n263_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n560_), .A2(new_n586_), .A3(new_n581_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n623_), .A2(new_n476_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(G29gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n373_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT43), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n534_), .A2(new_n535_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n623_), .B2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n432_), .A2(KEYINPUT43), .A3(new_n536_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n630_), .A2(new_n560_), .A3(new_n589_), .A4(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT44), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n432_), .A2(new_n536_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n559_), .B1(new_n635_), .B2(new_n628_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n636_), .A2(KEYINPUT44), .A3(new_n589_), .A4(new_n631_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n373_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT95), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(new_n639_), .A3(G29gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n638_), .B2(G29gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n627_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT96), .B(new_n627_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1328gat));
  NAND2_X1  g445(.A1(new_n634_), .A2(new_n637_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G36gat), .B1(new_n647_), .B2(new_n325_), .ZN(new_n648_));
  INV_X1    g447(.A(G36gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n625_), .A2(new_n649_), .A3(new_n597_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT45), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT46), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(G1329gat));
  NAND2_X1  g453(.A1(new_n606_), .A2(G43gat), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n625_), .A2(new_n606_), .ZN(new_n656_));
  OAI22_X1  g455(.A1(new_n647_), .A2(new_n655_), .B1(G43gat), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g457(.A1(new_n397_), .A2(G50gat), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT98), .Z(new_n660_));
  NAND2_X1  g459(.A1(new_n625_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n634_), .A2(new_n400_), .A3(new_n637_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT97), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n662_), .A2(new_n663_), .A3(G50gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n662_), .B2(G50gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(G1331gat));
  NAND2_X1  g465(.A1(new_n561_), .A2(new_n588_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT99), .Z(new_n668_));
  NOR2_X1   g467(.A1(new_n623_), .A2(new_n477_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT100), .Z(new_n671_));
  AOI21_X1  g470(.A(G57gat), .B1(new_n671_), .B2(new_n373_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n587_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n581_), .A2(new_n477_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR4_X1   g474(.A1(new_n623_), .A2(new_n560_), .A3(new_n673_), .A4(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(G57gat), .A3(new_n373_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT101), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n672_), .A2(new_n678_), .ZN(G1332gat));
  INV_X1    g478(.A(G64gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n671_), .A2(new_n680_), .A3(new_n597_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n676_), .B2(new_n597_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT48), .Z(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1333gat));
  NAND3_X1  g483(.A1(new_n671_), .A2(new_n233_), .A3(new_n606_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n676_), .A2(new_n606_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G71gat), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT102), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT102), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT49), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n688_), .A2(KEYINPUT49), .A3(new_n689_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n685_), .A2(new_n692_), .A3(new_n693_), .ZN(G1334gat));
  INV_X1    g493(.A(G78gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n671_), .A2(new_n695_), .A3(new_n400_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n676_), .A2(new_n400_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G78gat), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT103), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(KEYINPUT103), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n699_), .A2(KEYINPUT50), .A3(new_n700_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n696_), .A2(new_n703_), .A3(new_n704_), .ZN(G1335gat));
  NAND4_X1  g504(.A1(new_n669_), .A2(new_n560_), .A3(new_n586_), .A4(new_n588_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n496_), .A3(new_n373_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n630_), .A2(new_n560_), .A3(new_n631_), .A4(new_n674_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT105), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n373_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n712_), .B2(new_n496_), .ZN(G1336gat));
  AOI21_X1  g512(.A(G92gat), .B1(new_n708_), .B2(new_n597_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n597_), .A2(G92gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT106), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n711_), .B2(new_n716_), .ZN(G1337gat));
  OAI21_X1  g516(.A(G99gat), .B1(new_n710_), .B2(new_n263_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n706_), .B(KEYINPUT104), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n606_), .A2(new_n491_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n721_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT107), .B1(new_n708_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n718_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT51), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n718_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n708_), .A2(new_n492_), .A3(new_n400_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n629_), .B1(new_n423_), .B2(new_n431_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n560_), .B1(new_n732_), .B2(KEYINPUT43), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n628_), .B(new_n629_), .C1(new_n423_), .C2(new_n431_), .ZN(new_n734_));
  NOR4_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n397_), .A4(new_n675_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT108), .B1(new_n710_), .B2(new_n397_), .ZN(new_n738_));
  AND4_X1   g537(.A1(new_n731_), .A2(new_n737_), .A3(new_n738_), .A4(G106gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n492_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n731_), .B1(new_n740_), .B2(new_n738_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n730_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n730_), .B(new_n743_), .C1(new_n739_), .C2(new_n741_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1339gat));
  INV_X1    g546(.A(new_n586_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n477_), .A2(new_n578_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n562_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n567_), .A2(new_n750_), .A3(new_n569_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n570_), .A2(new_n562_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n570_), .A2(KEYINPUT55), .A3(new_n562_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT111), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n570_), .A2(new_n757_), .A3(KEYINPUT55), .A4(new_n562_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n759_), .A2(KEYINPUT113), .A3(KEYINPUT56), .A4(new_n575_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n759_), .A2(new_n575_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT112), .B(KEYINPUT56), .C1(new_n759_), .C2(new_n575_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n749_), .B1(new_n764_), .B2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n472_), .B1(new_n468_), .B2(new_n463_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT114), .B1(new_n462_), .B2(new_n466_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n464_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n462_), .A2(KEYINPUT114), .A3(new_n466_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n772_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n473_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT57), .B(new_n748_), .C1(new_n771_), .C2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n780_));
  AOI22_X1  g579(.A1(KEYINPUT111), .A2(new_n755_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n576_), .B1(new_n781_), .B2(new_n758_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT112), .B1(new_n782_), .B2(KEYINPUT56), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n766_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n783_), .A2(new_n784_), .A3(new_n762_), .A4(new_n763_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n476_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n778_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n780_), .B1(new_n787_), .B2(new_n586_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n779_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n776_), .A2(new_n473_), .A3(new_n578_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n766_), .A2(new_n767_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n760_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n536_), .B1(new_n792_), .B2(KEYINPUT58), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(KEYINPUT58), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT116), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n792_), .A2(KEYINPUT58), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n536_), .A4(new_n794_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n560_), .B1(new_n789_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n629_), .A2(new_n559_), .A3(new_n581_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n477_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n561_), .A2(new_n476_), .A3(new_n581_), .A4(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n801_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n373_), .ZN(new_n810_));
  NOR4_X1   g609(.A1(new_n597_), .A2(new_n810_), .A3(new_n400_), .A4(new_n263_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n793_), .A2(new_n795_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n560_), .B1(new_n789_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n808_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n811_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819_), .B2(new_n476_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n476_), .A2(G113gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n812_), .B2(new_n821_), .ZN(G1340gat));
  OAI21_X1  g621(.A(G120gat), .B1(new_n819_), .B2(new_n581_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n824_));
  AOI21_X1  g623(.A(G120gat), .B1(new_n588_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n824_), .B2(G120gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n809_), .A2(new_n811_), .A3(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT117), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n812_), .B2(new_n560_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n831_), .A2(KEYINPUT118), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(KEYINPUT118), .ZN(new_n833_));
  INV_X1    g632(.A(new_n819_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n560_), .A2(new_n830_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n832_), .A2(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1342gat));
  OAI21_X1  g635(.A(G134gat), .B1(new_n819_), .B2(new_n629_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n587_), .A2(G134gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n812_), .B2(new_n838_), .ZN(G1343gat));
  NOR2_X1   g638(.A1(new_n606_), .A2(new_n810_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n400_), .A3(new_n325_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n809_), .A2(KEYINPUT119), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n779_), .A2(new_n788_), .A3(new_n796_), .A4(new_n799_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n807_), .B1(new_n845_), .B2(new_n560_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n846_), .B2(new_n841_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n477_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT120), .B(G141gat), .Z(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n588_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT121), .B(G148gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n848_), .B2(new_n559_), .ZN(new_n858_));
  AOI211_X1 g657(.A(KEYINPUT122), .B(new_n560_), .C1(new_n843_), .C2(new_n847_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT119), .B1(new_n809_), .B2(new_n842_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n846_), .A2(new_n844_), .A3(new_n841_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n559_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT122), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n848_), .A2(new_n857_), .A3(new_n559_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n855_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n860_), .A2(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n848_), .A2(new_n868_), .A3(new_n673_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n629_), .B1(new_n843_), .B2(new_n847_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n868_), .ZN(G1347gat));
  NOR3_X1   g670(.A1(new_n325_), .A2(new_n400_), .A3(new_n425_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n816_), .A2(new_n477_), .A3(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(G169gat), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n816_), .A2(new_n872_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n476_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n874_), .A2(new_n876_), .B1(new_n281_), .B2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n874_), .B2(new_n876_), .ZN(G1348gat));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n809_), .A2(new_n881_), .A3(new_n397_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT124), .B1(new_n846_), .B2(new_n400_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n325_), .A2(new_n425_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n581_), .A2(new_n204_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n882_), .A2(new_n883_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n204_), .B1(new_n877_), .B2(new_n581_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT125), .ZN(G1349gat));
  NOR3_X1   g688(.A1(new_n877_), .A2(new_n285_), .A3(new_n560_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n882_), .A2(new_n883_), .A3(new_n559_), .A4(new_n884_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n220_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n877_), .B2(new_n629_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n673_), .A2(new_n222_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n877_), .B2(new_n894_), .ZN(G1351gat));
  NAND3_X1  g694(.A1(new_n398_), .A2(new_n263_), .A3(new_n597_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n846_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n477_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n588_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g700(.A1(new_n846_), .A2(new_n560_), .A3(new_n896_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT63), .B(G211gat), .Z(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n904_), .A2(KEYINPUT126), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(KEYINPUT126), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n902_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(G1354gat));
  AOI21_X1  g707(.A(G218gat), .B1(new_n897_), .B2(new_n673_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n536_), .A2(G218gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT127), .Z(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n897_), .B2(new_n911_), .ZN(G1355gat));
endmodule


