//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(G85gat), .B(G92gat), .Z(new_n204_));
  NOR2_X1   g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n204_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT8), .ZN(new_n212_));
  INV_X1    g011(.A(new_n210_), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  OR3_X1    g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT9), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n212_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(KEYINPUT11), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(G71gat), .ZN(new_n227_));
  INV_X1    g026(.A(G78gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n224_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n203_), .B1(new_n222_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT12), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n230_), .A2(new_n232_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n221_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n211_), .A2(KEYINPUT8), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n211_), .A2(KEYINPUT8), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n237_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n222_), .A2(new_n233_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT66), .A3(new_n237_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n240_), .A2(new_n249_), .A3(new_n241_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n221_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n238_), .A2(new_n237_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n245_), .A2(new_n247_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n236_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n203_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n246_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n222_), .A2(new_n233_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G120gat), .B(G148gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(G176gat), .B(G204gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n265_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n255_), .A2(new_n259_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(KEYINPUT13), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT13), .B1(new_n266_), .B2(new_n268_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n202_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n271_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(KEYINPUT69), .A3(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G29gat), .B(G36gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G43gat), .B(G50gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT15), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G15gat), .B(G22gat), .ZN(new_n280_));
  INV_X1    g079(.A(G1gat), .ZN(new_n281_));
  INV_X1    g080(.A(G8gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT14), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n280_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n283_), .A2(new_n284_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G8gat), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n279_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT75), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n289_), .A3(new_n278_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G229gat), .A2(G233gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n290_), .B(new_n278_), .Z(new_n296_));
  INV_X1    g095(.A(new_n294_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G113gat), .B(G141gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(G169gat), .B(G197gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n295_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT76), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n295_), .A2(new_n298_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n275_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G211gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(G218gat), .ZN(new_n309_));
  INV_X1    g108(.A(G218gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(G211gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT88), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(G211gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(G218gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n312_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n312_), .A2(new_n316_), .B1(new_n319_), .B2(new_n317_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT21), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n312_), .A2(new_n316_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n319_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT21), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT89), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT21), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n315_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n323_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n312_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n328_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT89), .B1(new_n333_), .B2(new_n324_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n327_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G141gat), .B(G148gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT84), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT84), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(G155gat), .A3(G162gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n338_), .B1(new_n343_), .B2(KEYINPUT1), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n337_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348_));
  INV_X1    g147(.A(G141gat), .ZN(new_n349_));
  INV_X1    g148(.A(G148gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n338_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n356_), .A2(new_n343_), .A3(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n347_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n336_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n335_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT90), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n359_), .A2(new_n360_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n321_), .A2(new_n325_), .ZN(new_n366_));
  OAI211_X1 g165(.A(G228gat), .B(G233gat), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT91), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT86), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n356_), .A2(new_n343_), .A3(new_n357_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n340_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n345_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n338_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n373_), .B1(new_n376_), .B2(new_n337_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n372_), .B1(new_n377_), .B2(KEYINPUT29), .ZN(new_n378_));
  INV_X1    g177(.A(new_n372_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n359_), .A2(new_n360_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT92), .ZN(new_n385_));
  INV_X1    g184(.A(new_n382_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n378_), .A2(new_n380_), .A3(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n383_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n384_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n370_), .A2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n364_), .B(new_n369_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  XOR2_X1   g195(.A(G127gat), .B(G134gat), .Z(new_n397_));
  INV_X1    g196(.A(G120gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G113gat), .ZN(new_n399_));
  INV_X1    g198(.A(G113gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G120gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G127gat), .B(G134gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G113gat), .B(G120gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n406_), .A3(KEYINPUT82), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n347_), .B2(new_n358_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n403_), .A2(new_n406_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n373_), .B(new_n412_), .C1(new_n376_), .C2(new_n337_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(KEYINPUT4), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT98), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT98), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n411_), .A2(new_n416_), .A3(new_n413_), .A4(KEYINPUT4), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n377_), .A2(new_n419_), .A3(new_n410_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT99), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n396_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(new_n218_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT0), .B(G57gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n411_), .A2(new_n413_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n396_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OR3_X1    g228(.A1(new_n422_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n426_), .B1(new_n422_), .B2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G183gat), .A2(G190gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT23), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT23), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G183gat), .A3(G190gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n435_), .A2(KEYINPUT80), .A3(G183gat), .A4(G190gat), .ZN(new_n439_));
  INV_X1    g238(.A(G190gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT77), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G190gat), .ZN(new_n443_));
  INV_X1    g242(.A(G183gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n438_), .A2(new_n439_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G169gat), .A2(G176gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT22), .ZN(new_n448_));
  AOI21_X1  g247(.A(G176gat), .B1(new_n448_), .B2(G169gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT78), .ZN(new_n450_));
  INV_X1    g249(.A(G169gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n448_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT79), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n449_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n453_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n455_), .B(KEYINPUT22), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n446_), .B(new_n447_), .C1(new_n456_), .C2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT25), .B(G183gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT26), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n463_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n462_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n434_), .A2(new_n436_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n447_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(G169gat), .A2(G176gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT24), .ZN(new_n470_));
  OR3_X1    g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n470_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n471_), .A4(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n461_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n461_), .A2(KEYINPUT81), .A3(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G71gat), .B(G99gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G43gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n478_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(new_n410_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G227gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(G15gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT30), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT31), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n482_), .A2(new_n487_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n432_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G64gat), .B(G92gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT96), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G8gat), .B(G36gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n496_), .B(KEYINPUT103), .Z(new_n497_));
  AOI21_X1  g296(.A(new_n326_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n333_), .A2(new_n324_), .A3(KEYINPUT89), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT20), .B1(new_n500_), .B2(new_n478_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT94), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n471_), .A2(new_n472_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G190gat), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n462_), .B2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n438_), .A2(new_n439_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n467_), .B1(G183gat), .B2(G190gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT22), .B(G169gat), .ZN(new_n508_));
  INV_X1    g307(.A(G176gat), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n468_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n505_), .A2(new_n506_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(new_n366_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n513_), .B(KEYINPUT20), .C1(new_n500_), .C2(new_n478_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n502_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n500_), .A2(new_n478_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n511_), .B2(new_n366_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n518_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n497_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT27), .ZN(new_n526_));
  INV_X1    g325(.A(new_n521_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n511_), .A2(new_n366_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(KEYINPUT20), .A3(new_n518_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n515_), .B2(new_n519_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n526_), .B1(new_n531_), .B2(new_n496_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n514_), .A2(new_n512_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n335_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n513_), .B1(new_n534_), .B2(KEYINPUT20), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n519_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n530_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n496_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n536_), .A2(KEYINPUT97), .A3(new_n496_), .A4(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n537_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n496_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n541_), .A3(new_n544_), .ZN(new_n545_));
  AOI221_X4 g344(.A(KEYINPUT104), .B1(new_n525_), .B2(new_n532_), .C1(new_n545_), .C2(new_n526_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT104), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n526_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n532_), .A2(new_n525_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n395_), .B(new_n490_), .C1(new_n546_), .C2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n488_), .A2(new_n489_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT83), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n418_), .A2(new_n421_), .A3(new_n396_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n431_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n431_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT101), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n431_), .A2(KEYINPUT101), .A3(new_n560_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n559_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n496_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n539_), .B2(new_n538_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n567_), .A3(new_n541_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n496_), .A2(KEYINPUT32), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n531_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n520_), .A2(new_n524_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n432_), .B(new_n570_), .C1(new_n571_), .C2(new_n569_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n394_), .B1(new_n568_), .B2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n392_), .A2(new_n430_), .A3(new_n393_), .A4(new_n431_), .ZN(new_n574_));
  AOI221_X4 g373(.A(new_n574_), .B1(new_n525_), .B2(new_n532_), .C1(new_n545_), .C2(new_n526_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n554_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n307_), .B1(new_n551_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT71), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT36), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n252_), .A2(new_n279_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n242_), .A2(new_n278_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n584_), .A2(KEYINPUT70), .A3(new_n585_), .A4(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n239_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n279_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT70), .B(new_n585_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n588_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n585_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT35), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n589_), .A2(new_n594_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT72), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n589_), .A2(new_n594_), .A3(new_n600_), .A4(new_n597_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n583_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n581_), .A2(KEYINPUT36), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n602_), .A2(KEYINPUT73), .B1(new_n603_), .B2(new_n598_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n582_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT73), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n604_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n598_), .A2(new_n583_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n598_), .A2(new_n603_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(KEYINPUT37), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n290_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n233_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT16), .ZN(new_n620_));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT17), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n618_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT17), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n618_), .B1(new_n625_), .B2(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n615_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n577_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n281_), .A3(new_n432_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT105), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n609_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n551_), .B2(new_n576_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n307_), .A2(new_n628_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n432_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G1gat), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n634_), .A2(new_n635_), .A3(new_n642_), .ZN(G1324gat));
  NOR2_X1   g442(.A1(new_n546_), .A2(new_n550_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n630_), .A2(new_n282_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(new_n644_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  AND4_X1   g446(.A1(KEYINPUT106), .A2(new_n646_), .A3(new_n647_), .A4(G8gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n282_), .B1(new_n649_), .B2(KEYINPUT39), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n646_), .A2(new_n650_), .B1(KEYINPUT106), .B2(new_n647_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n645_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g452(.A(new_n554_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n630_), .A2(new_n484_), .A3(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT107), .Z(new_n656_));
  OAI21_X1  g455(.A(G15gat), .B1(new_n640_), .B2(new_n554_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n657_), .A2(KEYINPUT41), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(KEYINPUT41), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n658_), .A3(new_n659_), .ZN(G1326gat));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n394_), .B(KEYINPUT108), .Z(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n639_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT42), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n630_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  NOR2_X1   g465(.A1(new_n609_), .A2(new_n627_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n577_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n432_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n275_), .A2(new_n628_), .A3(new_n306_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n551_), .A2(new_n576_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(KEYINPUT110), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(KEYINPUT110), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n674_), .A2(new_n615_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n614_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n681_), .B(new_n676_), .C1(new_n551_), .C2(new_n576_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n673_), .B1(new_n679_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n673_), .B(KEYINPUT44), .C1(new_n679_), .C2(new_n682_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n432_), .A2(G29gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n670_), .B1(new_n687_), .B2(new_n688_), .ZN(G1328gat));
  INV_X1    g488(.A(new_n644_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(G36gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n577_), .A2(new_n691_), .A3(new_n667_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT45), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n685_), .A2(new_n644_), .A3(new_n686_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n696_), .A2(new_n697_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n695_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1329gat));
  NAND4_X1  g501(.A1(new_n685_), .A2(G43gat), .A3(new_n552_), .A4(new_n686_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT112), .B(G43gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n668_), .B2(new_n554_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g506(.A(G50gat), .B1(new_n669_), .B2(new_n662_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n394_), .A2(G50gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n687_), .B2(new_n709_), .ZN(G1331gat));
  OR2_X1    g509(.A1(new_n275_), .A2(new_n306_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n576_), .B2(new_n551_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n629_), .ZN(new_n713_));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n432_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n711_), .A2(new_n628_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n637_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n641_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1332gat));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n713_), .A2(new_n720_), .A3(new_n644_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722_));
  INV_X1    g521(.A(new_n717_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n644_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(G64gat), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT48), .B(new_n720_), .C1(new_n723_), .C2(new_n644_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n721_), .B1(new_n725_), .B2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n654_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT113), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n713_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT49), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n723_), .A2(new_n654_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G71gat), .ZN(new_n734_));
  AOI211_X1 g533(.A(KEYINPUT49), .B(new_n728_), .C1(new_n723_), .C2(new_n654_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1334gat));
  NAND3_X1  g535(.A1(new_n713_), .A2(new_n228_), .A3(new_n662_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n723_), .A2(new_n662_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G78gat), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT50), .B(new_n228_), .C1(new_n723_), .C2(new_n662_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n711_), .A2(new_n627_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n679_), .B2(new_n682_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n641_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n712_), .A2(new_n667_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n218_), .A3(new_n432_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1336gat));
  OAI21_X1  g547(.A(G92gat), .B1(new_n744_), .B2(new_n690_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(new_n219_), .A3(new_n644_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1337gat));
  OAI21_X1  g550(.A(G99gat), .B1(new_n744_), .B2(new_n554_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n214_), .A3(new_n552_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n754_), .B(new_n755_), .Z(G1338gat));
  NAND3_X1  g555(.A1(new_n746_), .A2(new_n215_), .A3(new_n394_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n743_), .B(new_n394_), .C1(new_n679_), .C2(new_n682_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n215_), .B1(new_n759_), .B2(KEYINPUT52), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n758_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n758_), .B2(new_n761_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n757_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g564(.A(KEYINPUT58), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n252_), .A2(new_n253_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n258_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT66), .B1(new_n246_), .B2(new_n237_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n243_), .A2(new_n244_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n767_), .B(new_n768_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n256_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT118), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n774_), .A3(new_n256_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n767_), .B1(new_n770_), .B2(new_n769_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n234_), .B(KEYINPUT67), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n236_), .A2(new_n254_), .A3(KEYINPUT55), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n773_), .A2(new_n775_), .A3(new_n779_), .A4(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n265_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT121), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n265_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n265_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT121), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n292_), .A2(new_n293_), .A3(new_n297_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n301_), .B1(new_n296_), .B2(new_n294_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n303_), .A2(new_n268_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n789_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n766_), .B1(new_n785_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n793_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(KEYINPUT58), .C1(new_n784_), .C2(new_n783_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n798_), .A3(new_n615_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n266_), .A2(new_n268_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n303_), .A3(new_n792_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n268_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n781_), .B2(new_n265_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n805_), .B2(KEYINPUT56), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n804_), .B(new_n788_), .C1(new_n781_), .C2(new_n265_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n801_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n609_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT57), .B1(new_n808_), .B2(new_n609_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n799_), .B(new_n809_), .C1(new_n810_), .C2(KEYINPUT120), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n810_), .A2(KEYINPUT120), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n628_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n306_), .A2(new_n628_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n270_), .A2(new_n271_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n818_), .A2(KEYINPUT117), .A3(new_n819_), .A4(new_n681_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(new_n681_), .A3(new_n817_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(KEYINPUT54), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(KEYINPUT54), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n820_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n813_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n690_), .A2(new_n432_), .A3(new_n395_), .A4(new_n552_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT122), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n799_), .A2(new_n809_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n628_), .B1(new_n831_), .B2(new_n810_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n825_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n828_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(new_n306_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(G113gat), .ZN(new_n837_));
  INV_X1    g636(.A(new_n829_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(new_n400_), .A3(new_n306_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1340gat));
  INV_X1    g639(.A(new_n275_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n830_), .A2(new_n841_), .A3(new_n835_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n398_), .B1(new_n275_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n838_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n398_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1341gat));
  NAND3_X1  g645(.A1(new_n830_), .A2(new_n627_), .A3(new_n835_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G127gat), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n829_), .A2(G127gat), .A3(new_n628_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1342gat));
  NAND3_X1  g649(.A1(new_n830_), .A2(new_n615_), .A3(new_n835_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G134gat), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n829_), .A2(G134gat), .A3(new_n609_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1343gat));
  XNOR2_X1  g653(.A(KEYINPUT123), .B(G141gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n690_), .A2(new_n432_), .A3(new_n394_), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n654_), .B(new_n858_), .C1(new_n813_), .C2(new_n825_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n859_), .B2(new_n306_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n858_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n826_), .A2(new_n554_), .A3(new_n306_), .A4(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(KEYINPUT124), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n856_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n857_), .A3(new_n306_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(KEYINPUT124), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n855_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n859_), .A2(new_n841_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n859_), .A2(new_n627_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n859_), .B2(new_n636_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n615_), .A2(G162gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT125), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n859_), .B2(new_n876_), .ZN(G1347gat));
  AOI21_X1  g676(.A(new_n662_), .B1(new_n832_), .B2(new_n825_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n554_), .A2(new_n432_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n644_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n878_), .A2(new_n306_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n882_), .A2(new_n883_), .A3(new_n451_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n508_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n882_), .B2(new_n451_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(G1348gat));
  NAND3_X1  g686(.A1(new_n878_), .A2(new_n841_), .A3(new_n881_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n394_), .B1(new_n813_), .B2(new_n825_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n880_), .A2(new_n509_), .A3(new_n275_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n888_), .A2(new_n509_), .B1(new_n889_), .B2(new_n890_), .ZN(G1349gat));
  NOR2_X1   g690(.A1(new_n880_), .A2(new_n628_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G183gat), .B1(new_n889_), .B2(new_n892_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n880_), .A2(new_n628_), .A3(new_n462_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n878_), .B2(new_n894_), .ZN(G1350gat));
  NAND4_X1  g694(.A1(new_n878_), .A2(new_n636_), .A3(new_n504_), .A4(new_n881_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n878_), .A2(new_n615_), .A3(new_n881_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n440_), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n690_), .A2(new_n574_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n826_), .A2(new_n554_), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n306_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g701(.A1(new_n826_), .A2(new_n554_), .A3(new_n841_), .A4(new_n899_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(G204gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(KEYINPUT127), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n903_), .A2(new_n907_), .A3(G204gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n903_), .A2(new_n909_), .A3(G204gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n903_), .B2(G204gat), .ZN(new_n911_));
  OAI22_X1  g710(.A1(new_n906_), .A2(new_n908_), .B1(new_n910_), .B2(new_n911_), .ZN(G1353gat));
  NAND4_X1  g711(.A1(new_n826_), .A2(new_n627_), .A3(new_n554_), .A4(new_n899_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AND2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  NAND3_X1  g716(.A1(new_n900_), .A2(new_n310_), .A3(new_n636_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n900_), .A2(new_n615_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n310_), .ZN(G1355gat));
endmodule


