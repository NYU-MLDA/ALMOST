//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_;
  XNOR2_X1  g000(.A(KEYINPUT67), .B(G71gat), .ZN(new_n202_));
  INV_X1    g001(.A(G78gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT11), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n202_), .B(G78gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT66), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n217_), .A2(new_n220_), .A3(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT65), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  INV_X1    g030(.A(G92gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G85gat), .A2(G92gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n213_), .B1(new_n227_), .B2(new_n237_), .ZN(new_n238_));
  NOR4_X1   g037(.A1(new_n215_), .A2(new_n216_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n230_), .A2(new_n236_), .A3(new_n213_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n243_));
  INV_X1    g042(.A(G106gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT64), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n243_), .A2(new_n248_), .A3(new_n244_), .A4(new_n245_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT9), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n228_), .A2(new_n229_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(G85gat), .A3(G92gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n223_), .A2(new_n253_), .A3(new_n225_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n212_), .A2(new_n242_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n211_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G230gat), .ZN(new_n261_));
  INV_X1    g060(.A(G233gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT68), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n266_), .A3(new_n263_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n259_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n263_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n250_), .A2(KEYINPUT69), .A3(new_n255_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT69), .B1(new_n250_), .B2(new_n255_), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n271_), .A2(new_n272_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n268_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n269_), .A2(new_n270_), .A3(new_n257_), .A4(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n267_), .A3(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G120gat), .B(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT5), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G176gat), .B(G204gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n265_), .A2(new_n267_), .A3(new_n276_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT13), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT13), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G232gat), .A2(G233gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT34), .Z(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G43gat), .B(G50gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G43gat), .B(G50gat), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n293_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT15), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT15), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n256_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n250_), .A2(KEYINPUT69), .A3(new_n255_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n304_), .B1(new_n242_), .B2(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n256_), .B(new_n299_), .C1(new_n238_), .C2(new_n241_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n290_), .A2(new_n291_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n292_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n273_), .A2(new_n303_), .A3(new_n301_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n310_), .A2(new_n311_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n292_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G190gat), .B(G218gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(G134gat), .B(G162gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT36), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(KEYINPUT71), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n322_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT37), .ZN(new_n328_));
  INV_X1    g127(.A(new_n326_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n318_), .B(KEYINPUT71), .C1(new_n329_), .C2(new_n323_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n327_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n328_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G15gat), .B(G22gat), .ZN(new_n333_));
  INV_X1    g132(.A(G1gat), .ZN(new_n334_));
  INV_X1    g133(.A(G8gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT14), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G1gat), .B(G8gat), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n338_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G231gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(new_n211_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G127gat), .B(G155gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT16), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G183gat), .B(G211gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n349_), .B2(KEYINPUT17), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n344_), .A2(new_n350_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n349_), .A2(KEYINPUT17), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n331_), .A2(new_n332_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n288_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT73), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT1), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(G155gat), .A3(G162gat), .ZN(new_n362_));
  OR2_X1    g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G141gat), .B(G148gat), .Z(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(KEYINPUT2), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(KEYINPUT2), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT3), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n368_), .A2(new_n369_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n363_), .A2(new_n359_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n366_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n376_), .A2(KEYINPUT29), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT28), .Z(new_n378_));
  XOR2_X1   g177(.A(G22gat), .B(G50gat), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(KEYINPUT29), .ZN(new_n381_));
  INV_X1    g180(.A(G218gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G211gat), .ZN(new_n383_));
  INV_X1    g182(.A(G211gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G218gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n387_));
  INV_X1    g186(.A(G204gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT21), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(G197gat), .B2(G204gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n386_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(G197gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT84), .B(G197gat), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n391_), .B(new_n394_), .C1(new_n395_), .C2(new_n388_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n394_), .B1(new_n395_), .B2(new_n388_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT21), .A3(new_n386_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n381_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(G228gat), .A3(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n397_), .A2(new_n399_), .A3(KEYINPUT85), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n404_), .A2(new_n381_), .A3(new_n405_), .A4(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(KEYINPUT86), .Z(new_n409_));
  NAND3_X1  g208(.A1(new_n402_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n402_), .B2(new_n407_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n380_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n402_), .A2(new_n407_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n409_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n410_), .A3(new_n379_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n378_), .B1(new_n413_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n413_), .A2(new_n417_), .A3(new_n378_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G183gat), .A2(G190gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n427_));
  INV_X1    g226(.A(G169gat), .ZN(new_n428_));
  INV_X1    g227(.A(G176gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT24), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n426_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n430_), .A2(KEYINPUT24), .A3(new_n435_), .A4(new_n431_), .ZN(new_n436_));
  INV_X1    g235(.A(G183gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT25), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT25), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G183gat), .ZN(new_n440_));
  INV_X1    g239(.A(G190gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT26), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G190gat), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n438_), .A2(new_n440_), .A3(new_n442_), .A4(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n436_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n436_), .B2(new_n445_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n434_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n437_), .A2(new_n441_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n424_), .A2(new_n425_), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT22), .B(G169gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(KEYINPUT81), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT81), .B1(new_n428_), .B2(KEYINPUT22), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n429_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n435_), .B(new_n451_), .C1(new_n453_), .C2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n449_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G71gat), .B(G99gat), .ZN(new_n460_));
  INV_X1    g259(.A(G43gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G227gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(G15gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n462_), .B(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n449_), .A2(KEYINPUT30), .A3(new_n456_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n465_), .B1(new_n459_), .B2(new_n466_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT83), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n467_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G127gat), .B(G134gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G113gat), .B(G120gat), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OR3_X1    g277(.A1(new_n474_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n475_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT31), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n470_), .A2(new_n473_), .A3(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT83), .B(new_n482_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n421_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n457_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n489_));
  NAND2_X1  g288(.A1(G226gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n451_), .A2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n424_), .A2(new_n450_), .A3(KEYINPUT88), .A4(new_n425_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n452_), .A2(new_n429_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n493_), .A2(new_n435_), .A3(new_n494_), .A4(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n426_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n433_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n497_), .A2(new_n436_), .A3(new_n445_), .A4(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n400_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n491_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n488_), .A2(new_n503_), .A3(KEYINPUT20), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT89), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n397_), .A2(new_n399_), .A3(KEYINPUT85), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT85), .B1(new_n397_), .B2(new_n399_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n506_), .B1(new_n509_), .B2(new_n457_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n503_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n506_), .B1(new_n500_), .B2(new_n400_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n509_), .B2(new_n457_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n491_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G8gat), .B(G36gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(G64gat), .B(G92gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AND4_X1   g321(.A1(KEYINPUT91), .A2(new_n513_), .A3(new_n516_), .A4(new_n522_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n505_), .A2(new_n512_), .B1(new_n491_), .B2(new_n515_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n522_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT91), .B1(new_n524_), .B2(new_n522_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G1gat), .B(G29gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT0), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(G57gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(new_n231_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G225gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT92), .ZN(new_n534_));
  INV_X1    g333(.A(new_n376_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n481_), .B2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n479_), .A2(new_n480_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n537_), .A2(KEYINPUT92), .A3(new_n376_), .A4(new_n478_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n476_), .A2(new_n480_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(new_n376_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n536_), .A2(new_n538_), .A3(new_n541_), .A4(KEYINPUT4), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n481_), .A2(new_n535_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n533_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n533_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n540_), .B1(new_n543_), .B2(KEYINPUT92), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n547_), .B1(new_n548_), .B2(new_n536_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n532_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT33), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(KEYINPUT93), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n542_), .A2(new_n545_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n547_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n549_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(KEYINPUT93), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n532_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n553_), .B2(new_n547_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n542_), .A2(KEYINPUT94), .A3(new_n533_), .A4(new_n545_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n548_), .A2(new_n547_), .A3(new_n536_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n560_), .A2(new_n531_), .A3(new_n561_), .A4(new_n562_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n552_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n527_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n556_), .B(new_n532_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n500_), .B(KEYINPUT95), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n510_), .B1(new_n400_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n491_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n491_), .B2(new_n515_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n522_), .A2(KEYINPUT32), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n511_), .B1(new_n510_), .B2(new_n503_), .ZN(new_n573_));
  AND4_X1   g372(.A1(new_n511_), .A2(new_n488_), .A3(KEYINPUT20), .A4(new_n503_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n516_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n566_), .B(new_n572_), .C1(new_n575_), .C2(new_n571_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n487_), .B1(new_n565_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(new_n521_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT27), .A3(new_n525_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT96), .B1(new_n527_), .B2(KEYINPUT27), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n524_), .A2(KEYINPUT91), .A3(new_n522_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n575_), .B2(new_n521_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n575_), .A2(new_n521_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n582_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT96), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT27), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n580_), .B1(new_n581_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n420_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n485_), .B(new_n484_), .C1(new_n591_), .C2(new_n418_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n419_), .A2(new_n486_), .A3(new_n420_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n566_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n577_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT77), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n341_), .A2(new_n302_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n339_), .A2(new_n340_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n341_), .A2(new_n302_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n299_), .A2(new_n340_), .A3(new_n339_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(KEYINPUT74), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n602_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n301_), .A2(new_n303_), .A3(new_n341_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n601_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G169gat), .B(G197gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n613_), .A2(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n614_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n616_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n596_), .B1(new_n610_), .B2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n606_), .A2(new_n609_), .A3(KEYINPUT77), .A4(new_n622_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT78), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n610_), .B2(new_n623_), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT78), .B(new_n622_), .C1(new_n606_), .C2(new_n609_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n624_), .B(new_n625_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n358_), .A2(new_n595_), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n334_), .A3(new_n566_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT38), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n327_), .A2(KEYINPUT98), .A3(new_n330_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT98), .B1(new_n327_), .B2(new_n330_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n595_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n288_), .A2(new_n629_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n288_), .A2(KEYINPUT97), .A3(new_n629_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n355_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n638_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n566_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n633_), .A2(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649_));
  INV_X1    g448(.A(new_n590_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G8gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n652_), .B2(KEYINPUT39), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n651_), .A2(KEYINPUT99), .A3(new_n654_), .A4(G8gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(KEYINPUT39), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n653_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n631_), .A2(new_n335_), .A3(new_n650_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n486_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n644_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n631_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1326gat));
  INV_X1    g467(.A(G22gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n421_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n631_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n644_), .A2(new_n670_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(G22gat), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n669_), .B(new_n672_), .C1(new_n644_), .C2(new_n670_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n671_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT102), .Z(G1327gat));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n587_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n594_), .B(new_n579_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n565_), .A2(new_n576_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n487_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n331_), .A2(new_n332_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n680_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT43), .B(new_n688_), .C1(new_n683_), .C2(new_n686_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n641_), .A2(new_n642_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n355_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n679_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n595_), .B2(new_n688_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n687_), .A2(new_n680_), .A3(new_n689_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n698_), .A2(KEYINPUT44), .A3(new_n355_), .A4(new_n693_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n699_), .A3(new_n566_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G29gat), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n637_), .A2(new_n355_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n595_), .A2(new_n639_), .A3(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n646_), .A2(G29gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT103), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n706_), .ZN(G1328gat));
  NAND2_X1  g506(.A1(new_n695_), .A2(new_n699_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G36gat), .B1(new_n708_), .B2(new_n590_), .ZN(new_n709_));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n703_), .A2(new_n710_), .A3(new_n650_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT46), .Z(G1329gat));
  AOI21_X1  g513(.A(G43gat), .B1(new_n703_), .B2(new_n663_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n708_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n486_), .A2(new_n461_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g518(.A(G50gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n703_), .A2(new_n720_), .A3(new_n670_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(new_n670_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT104), .ZN(new_n723_));
  OAI21_X1  g522(.A(G50gat), .B1(new_n722_), .B2(KEYINPUT104), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n288_), .A2(new_n629_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n687_), .A2(new_n636_), .A3(new_n354_), .A4(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT106), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(G57gat), .A3(new_n566_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT107), .Z(new_n730_));
  INV_X1    g529(.A(new_n288_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n356_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n630_), .B1(new_n732_), .B2(KEYINPUT105), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n595_), .B(new_n733_), .C1(KEYINPUT105), .C2(new_n732_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n566_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n730_), .A2(new_n735_), .ZN(G1332gat));
  INV_X1    g535(.A(G64gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n728_), .B2(new_n650_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n739_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n734_), .A2(new_n737_), .A3(new_n650_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n740_), .A2(new_n741_), .A3(new_n742_), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n728_), .B2(new_n663_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n486_), .A2(G71gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT110), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n734_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1334gat));
  AOI21_X1  g550(.A(new_n203_), .B1(new_n728_), .B2(new_n670_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n734_), .A2(new_n203_), .A3(new_n670_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1335gat));
  NOR4_X1   g555(.A1(new_n595_), .A2(new_n629_), .A3(new_n288_), .A4(new_n702_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n231_), .A3(new_n566_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n726_), .A2(new_n355_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT112), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n760_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n646_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n758_), .B1(new_n765_), .B2(new_n231_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n757_), .A2(new_n232_), .A3(new_n650_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n590_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n232_), .ZN(G1337gat));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n763_), .B1(new_n698_), .B2(new_n760_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n764_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n663_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G99gat), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n243_), .A2(new_n245_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n757_), .A2(new_n663_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT113), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n486_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n778_));
  INV_X1    g577(.A(G99gat), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT113), .B(new_n776_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n770_), .B(KEYINPUT51), .C1(new_n777_), .C2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n786_), .B2(new_n780_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n784_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT114), .B1(new_n788_), .B2(new_n783_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n782_), .B1(new_n787_), .B2(new_n789_), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n757_), .A2(new_n244_), .A3(new_n670_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  INV_X1    g591(.A(new_n761_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n670_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n794_), .B2(G106gat), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT52), .B(new_n244_), .C1(new_n793_), .C2(new_n670_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g597(.A1(new_n592_), .A2(new_n646_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n629_), .A2(new_n284_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n276_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n269_), .A2(new_n257_), .A3(new_n275_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n263_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n802_), .B1(new_n276_), .B2(new_n801_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n281_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT56), .B(new_n281_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n800_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n610_), .A2(new_n623_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT78), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n610_), .A2(new_n626_), .A3(new_n623_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n608_), .B(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n602_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n602_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n623_), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n814_), .A2(new_n815_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n285_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n636_), .B(KEYINPUT57), .C1(new_n812_), .C2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT117), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n629_), .A2(new_n284_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n811_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n276_), .A2(new_n801_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT55), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n281_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n825_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n285_), .A2(new_n821_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(KEYINPUT57), .A4(new_n636_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n824_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n821_), .A2(new_n284_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n838_), .A2(KEYINPUT58), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n688_), .B1(new_n838_), .B2(KEYINPUT58), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n636_), .B1(new_n812_), .B2(new_n822_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n839_), .A2(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n354_), .B1(new_n836_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n288_), .A2(new_n630_), .A3(new_n356_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n590_), .B(new_n799_), .C1(new_n844_), .C2(new_n847_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n848_), .A2(KEYINPUT118), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(KEYINPUT118), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n629_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT119), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n848_), .A2(new_n857_), .A3(KEYINPUT59), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n854_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n629_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n853_), .B1(new_n861_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n859_), .B2(new_n731_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n731_), .A2(new_n865_), .A3(new_n863_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n865_), .B2(new_n863_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n849_), .A2(new_n850_), .A3(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT120), .B1(new_n864_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n854_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n858_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n857_), .B1(new_n848_), .B2(KEYINPUT59), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n870_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G120gat), .B1(new_n873_), .B2(new_n288_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875_));
  INV_X1    g674(.A(new_n868_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n869_), .A2(new_n877_), .ZN(G1341gat));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n851_), .A2(new_n879_), .A3(new_n354_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n859_), .A2(new_n354_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n882_), .B2(new_n879_), .ZN(G1342gat));
  INV_X1    g682(.A(G134gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n851_), .A2(new_n884_), .A3(new_n637_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n859_), .A2(new_n689_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n887_), .B2(new_n884_), .ZN(G1343gat));
  OR2_X1    g687(.A1(new_n844_), .A2(new_n847_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n889_), .A2(new_n590_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n646_), .A2(new_n593_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n630_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT121), .B(G141gat), .Z(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n288_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g696(.A1(new_n892_), .A2(new_n355_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G155gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n892_), .B2(new_n688_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n636_), .A2(G162gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n892_), .B2(new_n902_), .ZN(G1347gat));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n590_), .A2(new_n566_), .A3(new_n592_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n629_), .B(new_n905_), .C1(new_n844_), .C2(new_n847_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT122), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n889_), .A2(new_n905_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n452_), .A3(new_n629_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(KEYINPUT62), .B1(new_n907_), .B2(G169gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n904_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n912_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n914_), .A2(KEYINPUT123), .A3(new_n908_), .A4(new_n910_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1348gat));
  NAND2_X1  g715(.A1(new_n909_), .A2(new_n731_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g717(.A1(new_n909_), .A2(new_n354_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G183gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n438_), .A2(new_n440_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n919_), .ZN(G1350gat));
  AOI21_X1  g721(.A(new_n441_), .B1(new_n909_), .B2(new_n689_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT124), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n909_), .A2(new_n442_), .A3(new_n444_), .A4(new_n637_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n844_), .A2(new_n847_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n593_), .A2(new_n566_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT125), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n927_), .A2(new_n590_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n629_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n731_), .ZN(new_n933_));
  XOR2_X1   g732(.A(KEYINPUT126), .B(G204gat), .Z(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1353gat));
  NAND2_X1  g734(.A1(new_n930_), .A2(new_n354_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT63), .B(G211gat), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(KEYINPUT127), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n936_), .A2(new_n940_), .A3(new_n937_), .ZN(new_n941_));
  AOI211_X1 g740(.A(KEYINPUT63), .B(G211gat), .C1(new_n930_), .C2(new_n354_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n939_), .A2(new_n941_), .A3(new_n942_), .ZN(G1354gat));
  NAND3_X1  g742(.A1(new_n930_), .A2(new_n382_), .A3(new_n637_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n930_), .A2(new_n689_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n944_), .B1(new_n946_), .B2(new_n382_), .ZN(G1355gat));
endmodule


