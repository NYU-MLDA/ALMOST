//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n203_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT79), .B1(new_n212_), .B2(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(new_n213_), .C1(new_n214_), .C2(KEYINPUT79), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(G169gat), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n210_), .A2(new_n215_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT30), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G15gat), .B(G43gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT31), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n222_), .A2(new_n223_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G227gat), .A2(G233gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(G71gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G99gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G127gat), .B(G134gat), .Z(new_n232_));
  XOR2_X1   g031(.A(G113gat), .B(G120gat), .Z(new_n233_));
  XOR2_X1   g032(.A(new_n232_), .B(new_n233_), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n231_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OR3_X1    g035(.A1(new_n225_), .A2(new_n226_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242_));
  INV_X1    g041(.A(G155gat), .ZN(new_n243_));
  INV_X1    g042(.A(G162gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G155gat), .A2(G162gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n252_));
  INV_X1    g051(.A(G141gat), .ZN(new_n253_));
  INV_X1    g052(.A(G148gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT84), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n253_), .B(new_n254_), .C1(new_n255_), .C2(KEYINPUT3), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n257_), .B(KEYINPUT84), .C1(G141gat), .C2(G148gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n253_), .A2(new_n254_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT2), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n252_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n263_), .B(KEYINPUT85), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n256_), .A2(new_n258_), .B1(new_n260_), .B2(KEYINPUT2), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT86), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n251_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n247_), .B1(new_n272_), .B2(new_n249_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n248_), .A2(KEYINPUT1), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  AOI211_X1 g075(.A(new_n260_), .B(new_n271_), .C1(new_n273_), .C2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n234_), .B1(new_n270_), .B2(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT86), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT86), .B1(new_n267_), .B2(new_n268_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n250_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n234_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n273_), .A2(new_n276_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n260_), .A2(new_n271_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n282_), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n278_), .A2(new_n286_), .A3(KEYINPUT4), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n285_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n234_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n241_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G29gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(G85gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT0), .B(G57gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  NAND2_X1  g094(.A1(new_n278_), .A2(new_n286_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n296_), .A2(new_n241_), .ZN(new_n297_));
  OR3_X1    g096(.A1(new_n291_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n291_), .B2(new_n297_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n240_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT88), .ZN(new_n303_));
  INV_X1    g102(.A(G204gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(G197gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G197gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n306_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G218gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G211gat), .ZN(new_n318_));
  INV_X1    g117(.A(G211gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G218gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT89), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT21), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n316_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT21), .B1(new_n311_), .B2(new_n315_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n307_), .A2(new_n310_), .A3(new_n308_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT21), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(G197gat), .B2(G204gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n324_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n323_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n328_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n305_), .B1(new_n314_), .B2(G197gat), .ZN(new_n338_));
  NOR4_X1   g137(.A1(new_n312_), .A2(new_n313_), .A3(new_n303_), .A4(new_n310_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n330_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n322_), .A2(new_n324_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT90), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n327_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT29), .B1(new_n270_), .B2(new_n277_), .ZN(new_n344_));
  INV_X1    g143(.A(G228gat), .ZN(new_n345_));
  INV_X1    g144(.A(G233gat), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n343_), .B(new_n344_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT91), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n288_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n343_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT92), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n345_), .A2(new_n346_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n347_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G78gat), .B(G106gat), .Z(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n357_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n359_), .B(new_n347_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n288_), .A2(KEYINPUT29), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G22gat), .B(G50gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n358_), .A2(new_n366_), .A3(new_n360_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n327_), .B(new_n219_), .C1(new_n337_), .C2(new_n342_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT94), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT20), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n218_), .B(KEYINPUT97), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n216_), .ZN(new_n378_));
  XOR2_X1   g177(.A(KEYINPUT26), .B(G190gat), .Z(new_n379_));
  INV_X1    g178(.A(KEYINPUT95), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n214_), .A2(KEYINPUT95), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n211_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n210_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(KEYINPUT96), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT96), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n383_), .B2(new_n210_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n378_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n343_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n376_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n375_), .B1(new_n374_), .B2(KEYINPUT20), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n373_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT18), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n394_), .B(new_n395_), .Z(new_n396_));
  INV_X1    g195(.A(new_n373_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n388_), .B2(new_n343_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n336_), .B1(new_n328_), .B2(new_n335_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n340_), .A2(KEYINPUT90), .A3(new_n341_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n326_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT20), .B1(new_n401_), .B2(new_n219_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n392_), .A2(new_n396_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT98), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n392_), .A2(KEYINPUT98), .A3(new_n396_), .A4(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n392_), .A2(new_n403_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n396_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n404_), .A2(KEYINPUT27), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n401_), .B2(new_n219_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n416_), .A2(new_n375_), .B1(new_n343_), .B2(new_n388_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n391_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n397_), .A3(new_n418_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n401_), .A2(new_n378_), .A3(new_n384_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n373_), .B1(new_n420_), .B2(new_n402_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n409_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n414_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n413_), .A2(new_n424_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n302_), .A2(new_n370_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n300_), .B1(new_n414_), .B2(new_n423_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n358_), .A2(new_n366_), .A3(new_n360_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n366_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n413_), .B(new_n427_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n370_), .A2(KEYINPUT102), .A3(new_n413_), .A4(new_n427_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n287_), .A2(new_n290_), .A3(new_n241_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n295_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n296_), .A2(KEYINPUT99), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n241_), .B1(new_n296_), .B2(KEYINPUT99), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n299_), .A2(KEYINPUT33), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n441_), .B(new_n295_), .C1(new_n291_), .C2(new_n297_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n439_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n443_), .A2(new_n407_), .A3(new_n410_), .A4(new_n406_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n396_), .A2(KEYINPUT32), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n422_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT101), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT101), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n422_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n300_), .A3(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n398_), .A2(new_n402_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n417_), .A2(new_n418_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n452_), .B1(new_n453_), .B2(new_n373_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT100), .B1(new_n454_), .B2(new_n445_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT100), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n408_), .A2(new_n456_), .A3(new_n446_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n444_), .B1(new_n451_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n428_), .A2(new_n429_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n432_), .A2(new_n433_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n426_), .B1(new_n462_), .B2(new_n239_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G169gat), .B(G197gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G15gat), .B(G22gat), .Z(new_n468_));
  NAND2_X1  g267(.A1(G1gat), .A2(G8gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(KEYINPUT14), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT76), .ZN(new_n471_));
  XOR2_X1   g270(.A(G1gat), .B(G8gat), .Z(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n471_), .B(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G29gat), .B(G36gat), .Z(new_n475_));
  XOR2_X1   g274(.A(G43gat), .B(G50gat), .Z(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n471_), .B(new_n472_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n477_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n471_), .A2(new_n472_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n471_), .A2(new_n472_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n485_), .B1(new_n491_), .B2(new_n479_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n467_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT78), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n480_), .A2(new_n477_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n486_), .B1(new_n495_), .B2(new_n490_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(new_n466_), .C1(new_n484_), .C2(new_n486_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT78), .B(new_n467_), .C1(new_n487_), .C2(new_n492_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n463_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G85gat), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT66), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(KEYINPUT66), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT6), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(G99gat), .A3(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT10), .B(G99gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(G106gat), .ZN(new_n520_));
  OR3_X1    g319(.A1(new_n512_), .A2(new_n513_), .A3(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n513_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n505_), .A2(KEYINPUT68), .A3(new_n507_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT67), .ZN(new_n525_));
  NOR3_X1   g324(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n523_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI211_X1 g329(.A(KEYINPUT8), .B(new_n523_), .C1(new_n525_), .C2(new_n527_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n521_), .B(new_n522_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n482_), .A2(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n512_), .A2(new_n520_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n478_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G232gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT34), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT35), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n533_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(KEYINPUT35), .A3(new_n538_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(KEYINPUT36), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n538_), .A2(KEYINPUT35), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n533_), .A2(new_n536_), .A3(new_n546_), .A4(new_n539_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n541_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n544_), .B(KEYINPUT36), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n541_), .B2(new_n547_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT75), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT37), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT77), .B1(new_n562_), .B2(KEYINPUT17), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(new_n474_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT69), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n568_), .B2(KEYINPUT11), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(G57gat), .B(G64gat), .Z(new_n572_));
  INV_X1    g371(.A(KEYINPUT11), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n567_), .A3(KEYINPUT11), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n570_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n568_), .A2(new_n567_), .A3(KEYINPUT11), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n568_), .A2(KEYINPUT11), .ZN(new_n578_));
  OAI22_X1  g377(.A1(new_n577_), .A2(new_n569_), .B1(new_n578_), .B2(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n566_), .A2(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n562_), .A2(KEYINPUT17), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n566_), .A2(new_n580_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n558_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n535_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n580_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n580_), .A2(new_n591_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n590_), .A2(new_n591_), .B1(new_n532_), .B2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n580_), .B(new_n535_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n594_), .A2(KEYINPUT73), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT73), .B1(new_n594_), .B2(new_n598_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n593_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n534_), .A2(new_n602_), .A3(new_n535_), .A4(new_n580_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n594_), .A2(KEYINPUT70), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n590_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n597_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n606_), .A2(KEYINPUT71), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(KEYINPUT71), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n601_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT5), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n601_), .B(new_n615_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT13), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(KEYINPUT13), .A3(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n587_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n502_), .A2(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n623_), .A2(G1gat), .A3(new_n301_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n463_), .B2(new_n552_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n552_), .ZN(new_n629_));
  AOI22_X1  g428(.A1(new_n430_), .A2(new_n431_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n240_), .B1(new_n630_), .B2(new_n433_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT104), .B(new_n629_), .C1(new_n631_), .C2(new_n426_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n585_), .B1(new_n628_), .B2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n621_), .A2(new_n501_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n300_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(G1gat), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n626_), .A2(new_n636_), .ZN(G1324gat));
  XNOR2_X1  g436(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n628_), .A2(new_n632_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n425_), .A3(new_n584_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT106), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G8gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n641_), .B1(new_n628_), .B2(new_n632_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT106), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n646_), .A3(KEYINPUT39), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n648_));
  INV_X1    g447(.A(new_n425_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(G8gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n623_), .B2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n502_), .A2(KEYINPUT105), .A3(new_n622_), .A4(new_n650_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n647_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT39), .B1(new_n642_), .B2(new_n646_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n639_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n642_), .A2(new_n646_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n660_), .A2(new_n647_), .A3(new_n654_), .A4(new_n638_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n661_), .ZN(G1325gat));
  OR3_X1    g461(.A1(new_n623_), .A2(G15gat), .A3(new_n239_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n628_), .A2(new_n632_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n664_), .A2(new_n634_), .A3(new_n240_), .A4(new_n584_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n665_), .B2(G15gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT108), .B(new_n663_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1326gat));
  OR3_X1    g471(.A1(new_n623_), .A2(G22gat), .A3(new_n460_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n633_), .A2(new_n634_), .A3(new_n370_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(G22gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1327gat));
  NOR3_X1   g477(.A1(new_n621_), .A2(new_n629_), .A3(new_n584_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n502_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n300_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n558_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n463_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n685_), .B(new_n558_), .C1(new_n631_), .C2(new_n426_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n634_), .A2(new_n585_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n691_), .B(new_n688_), .C1(new_n684_), .C2(new_n686_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n300_), .A2(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n682_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  NOR2_X1   g494(.A1(new_n649_), .A2(G36gat), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OR3_X1    g496(.A1(new_n680_), .A2(KEYINPUT45), .A3(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT45), .B1(new_n680_), .B2(new_n697_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n690_), .A2(new_n692_), .A3(new_n649_), .ZN(new_n701_));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(KEYINPUT46), .B(new_n700_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  AND2_X1   g506(.A1(new_n240_), .A2(G43gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n693_), .A2(new_n708_), .ZN(new_n709_));
  XOR2_X1   g508(.A(KEYINPUT109), .B(G43gat), .Z(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n680_), .B2(new_n239_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(new_n715_), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1330gat));
  AOI21_X1  g516(.A(G50gat), .B1(new_n681_), .B2(new_n370_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n370_), .A2(G50gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n693_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(new_n621_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n500_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n633_), .A2(new_n300_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G57gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n463_), .A2(new_n500_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n621_), .A3(new_n586_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n301_), .A2(G57gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n726_), .B2(new_n727_), .ZN(G1332gat));
  OR3_X1    g527(.A1(new_n726_), .A2(G64gat), .A3(new_n649_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n633_), .A2(new_n425_), .A3(new_n722_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(G64gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n730_), .B2(G64gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(G1333gat));
  OR3_X1    g533(.A1(new_n726_), .A2(G71gat), .A3(new_n239_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n664_), .A2(new_n240_), .A3(new_n584_), .A4(new_n722_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G71gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT110), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n735_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1334gat));
  OR3_X1    g543(.A1(new_n726_), .A2(G78gat), .A3(new_n460_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n633_), .A2(new_n370_), .A3(new_n722_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G78gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G78gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1335gat));
  NOR3_X1   g549(.A1(new_n721_), .A2(new_n629_), .A3(new_n584_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n725_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n503_), .B1(new_n752_), .B2(new_n301_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT111), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n722_), .A2(new_n585_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n757_), .A2(new_n503_), .A3(new_n301_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n754_), .A2(new_n758_), .ZN(G1336gat));
  OAI21_X1  g558(.A(G92gat), .B1(new_n757_), .B2(new_n649_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n752_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n504_), .A3(new_n425_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1337gat));
  NAND2_X1  g562(.A1(new_n756_), .A2(new_n240_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G99gat), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n752_), .A2(new_n519_), .A3(new_n239_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT113), .ZN(new_n770_));
  INV_X1    g569(.A(G99gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n756_), .B2(new_n240_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n767_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n766_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n773_), .B2(new_n766_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT112), .B(KEYINPUT51), .C1(new_n772_), .C2(new_n767_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n776_), .A2(new_n780_), .ZN(G1338gat));
  INV_X1    g580(.A(G106gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n761_), .A2(new_n782_), .A3(new_n370_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n756_), .A2(new_n370_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(G106gat), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT52), .B(new_n782_), .C1(new_n756_), .C2(new_n370_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n783_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  NAND2_X1  g591(.A1(new_n500_), .A2(G113gat), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n601_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT115), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n601_), .A2(new_n797_), .A3(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n593_), .B(KEYINPUT55), .C1(new_n599_), .C2(new_n600_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n590_), .A2(new_n591_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n532_), .A2(new_n592_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n801_), .A2(new_n603_), .A3(new_n802_), .A4(new_n604_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n803_), .A2(KEYINPUT116), .A3(new_n597_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT116), .B1(new_n803_), .B2(new_n597_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n800_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n613_), .B1(new_n799_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT56), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n613_), .C1(new_n799_), .C2(new_n806_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n808_), .A2(new_n616_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n485_), .B1(new_n495_), .B2(new_n490_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n467_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n485_), .B1(new_n484_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n479_), .A2(new_n483_), .A3(KEYINPUT117), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n814_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n497_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n812_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n816_), .A2(new_n817_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT118), .B(new_n497_), .C1(new_n821_), .C2(new_n814_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n811_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n823_), .A2(new_n808_), .A3(new_n616_), .A4(new_n810_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n683_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n824_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n808_), .A2(new_n500_), .A3(new_n616_), .A4(new_n810_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n823_), .A2(new_n617_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n629_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(KEYINPUT57), .A3(new_n629_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n830_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n585_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n586_), .A2(new_n501_), .A3(new_n620_), .A4(new_n619_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n841_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n721_), .A2(new_n501_), .A3(new_n586_), .A4(new_n843_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n842_), .A2(new_n844_), .B1(KEYINPUT114), .B2(KEYINPUT54), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n839_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n649_), .A2(new_n300_), .A3(new_n460_), .A4(new_n240_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT120), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n849_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n793_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G113gat), .B1(new_n850_), .B2(new_n500_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n856_), .A2(KEYINPUT121), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(KEYINPUT121), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n855_), .B1(new_n857_), .B2(new_n858_), .ZN(G1340gat));
  XNOR2_X1  g658(.A(new_n852_), .B(KEYINPUT59), .ZN(new_n860_));
  OAI21_X1  g659(.A(G120gat), .B1(new_n860_), .B2(new_n721_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n721_), .A2(KEYINPUT60), .ZN(new_n862_));
  MUX2_X1   g661(.A(new_n862_), .B(KEYINPUT60), .S(G120gat), .Z(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT122), .B1(new_n850_), .B2(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n850_), .A2(KEYINPUT122), .A3(new_n863_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n861_), .B1(new_n864_), .B2(new_n865_), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n860_), .B2(new_n585_), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n852_), .A2(G127gat), .A3(new_n585_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1342gat));
  OAI21_X1  g668(.A(G134gat), .B1(new_n860_), .B2(new_n683_), .ZN(new_n870_));
  OR3_X1    g669(.A1(new_n852_), .A2(G134gat), .A3(new_n629_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1343gat));
  NOR3_X1   g671(.A1(new_n425_), .A2(new_n301_), .A3(new_n240_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n833_), .B2(new_n629_), .ZN(new_n874_));
  AOI211_X1 g673(.A(new_n835_), .B(new_n552_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n584_), .B1(new_n876_), .B2(new_n830_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n370_), .B(new_n873_), .C1(new_n877_), .C2(new_n845_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT123), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n847_), .A2(new_n880_), .A3(new_n370_), .A4(new_n873_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n500_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n621_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n584_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  AOI211_X1 g688(.A(new_n244_), .B(new_n683_), .C1(new_n879_), .C2(new_n881_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n882_), .A2(new_n552_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(KEYINPUT124), .A3(new_n244_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n629_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(G162gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n890_), .B1(new_n892_), .B2(new_n895_), .ZN(G1347gat));
  NOR3_X1   g695(.A1(new_n649_), .A2(new_n302_), .A3(new_n370_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n847_), .A2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT125), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT22), .B(G169gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n500_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n898_), .ZN(new_n902_));
  AOI211_X1 g701(.A(KEYINPUT62), .B(new_n204_), .C1(new_n902_), .C2(new_n500_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n500_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(G169gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n901_), .B1(new_n903_), .B2(new_n906_), .ZN(G1348gat));
  OAI21_X1  g706(.A(G176gat), .B1(new_n898_), .B2(new_n721_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n898_), .B(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n621_), .A2(new_n205_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n908_), .B1(new_n910_), .B2(new_n911_), .ZN(G1349gat));
  AOI21_X1  g711(.A(G183gat), .B1(new_n902_), .B2(new_n584_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n585_), .A2(new_n211_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n899_), .B2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n910_), .B2(new_n683_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n552_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n910_), .B2(new_n917_), .ZN(G1351gat));
  XNOR2_X1  g717(.A(KEYINPUT126), .B(G197gat), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n310_), .A2(KEYINPUT126), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n460_), .B1(new_n839_), .B2(new_n846_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n649_), .A2(new_n300_), .A3(new_n240_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n501_), .ZN(new_n924_));
  MUX2_X1   g723(.A(new_n919_), .B(new_n920_), .S(new_n924_), .Z(G1352gat));
  OAI21_X1  g724(.A(new_n304_), .B1(new_n923_), .B2(new_n721_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n921_), .A2(new_n621_), .A3(new_n309_), .A4(new_n922_), .ZN(new_n928_));
  AND3_X1   g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1353gat));
  NOR2_X1   g730(.A1(new_n923_), .A2(new_n585_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n932_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n933_));
  XOR2_X1   g732(.A(KEYINPUT63), .B(G211gat), .Z(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n932_), .B2(new_n934_), .ZN(G1354gat));
  OAI21_X1  g734(.A(G218gat), .B1(new_n923_), .B2(new_n683_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n552_), .A2(new_n317_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n923_), .B2(new_n937_), .ZN(G1355gat));
endmodule


