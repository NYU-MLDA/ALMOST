//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_,
    new_n983_, new_n984_;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT88), .B(G43gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n204_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT89), .B(G15gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n206_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n205_), .A2(new_n207_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n206_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n210_), .B1(new_n216_), .B2(new_n208_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n202_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT30), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT83), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT83), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G169gat), .A3(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(KEYINPUT22), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT22), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT86), .A3(G169gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n229_), .A2(G169gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(KEYINPUT85), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n225_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n225_), .B(KEYINPUT87), .C1(new_n235_), .C2(new_n232_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT23), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(G183gat), .B2(G190gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT26), .B(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(G183gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT25), .B1(new_n245_), .B2(KEYINPUT82), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(G183gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n244_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n252_), .A2(new_n221_), .A3(new_n223_), .A4(KEYINPUT24), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT84), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT84), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n252_), .A2(KEYINPUT24), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(new_n241_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n219_), .B1(new_n243_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n211_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n216_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT90), .A3(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n243_), .A2(new_n260_), .A3(new_n219_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n218_), .A2(new_n262_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT90), .B1(new_n263_), .B2(new_n264_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n266_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(new_n261_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(KEYINPUT91), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT31), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G113gat), .B(G120gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n267_), .A2(new_n270_), .A3(KEYINPUT91), .A4(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n272_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n275_), .B1(new_n272_), .B2(new_n277_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G141gat), .A2(G148gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(KEYINPUT1), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n286_), .B1(new_n288_), .B2(KEYINPUT1), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT92), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n287_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(G155gat), .B2(G162gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(KEYINPUT92), .A3(new_n286_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n285_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n286_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(new_n288_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n281_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n297_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT29), .B1(new_n295_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G228gat), .A2(G233gat), .ZN(new_n308_));
  INV_X1    g107(.A(G197gat), .ZN(new_n309_));
  INV_X1    g108(.A(G204gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G197gat), .A2(G204gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT21), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(KEYINPUT21), .A3(new_n312_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n316_), .A2(new_n317_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT93), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n307_), .A2(new_n308_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n308_), .B1(new_n307_), .B2(new_n320_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G78gat), .B(G106gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT94), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n324_), .A2(KEYINPUT97), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n321_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G22gat), .B(G50gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n330_));
  INV_X1    g129(.A(G155gat), .ZN(new_n331_));
  INV_X1    g130(.A(G162gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT1), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n290_), .B1(new_n333_), .B2(new_n296_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n287_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n294_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n300_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n337_), .A2(new_n303_), .A3(new_n304_), .A4(new_n298_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n297_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n336_), .A2(new_n284_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n330_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NOR4_X1   g141(.A1(new_n295_), .A2(new_n306_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n329_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(new_n339_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n293_), .A2(KEYINPUT92), .A3(new_n286_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT92), .B1(new_n293_), .B2(new_n286_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n287_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n341_), .B(new_n345_), .C1(new_n348_), .C2(new_n285_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT28), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n330_), .A3(new_n341_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n328_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n344_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n327_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n308_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n336_), .A2(new_n284_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n341_), .B1(new_n356_), .B2(new_n345_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n320_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n355_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n307_), .A2(new_n308_), .A3(new_n320_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n326_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n354_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT96), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n324_), .A2(KEYINPUT95), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n361_), .A2(new_n365_), .B1(new_n344_), .B2(new_n352_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n324_), .A2(KEYINPUT95), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n359_), .A2(new_n360_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n364_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n365_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n371_));
  AND4_X1   g170(.A1(new_n364_), .A2(new_n353_), .A3(new_n371_), .A4(new_n369_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n363_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT98), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n353_), .A2(new_n371_), .A3(new_n369_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT96), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n353_), .A2(new_n371_), .A3(new_n364_), .A4(new_n369_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT98), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(new_n363_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n275_), .B1(new_n295_), .B2(new_n306_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n273_), .B(new_n274_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n345_), .B(new_n383_), .C1(new_n348_), .C2(new_n285_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n384_), .A3(KEYINPUT4), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT104), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT104), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n382_), .A2(new_n384_), .A3(new_n391_), .A4(KEYINPUT4), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n275_), .B(new_n393_), .C1(new_n295_), .C2(new_n306_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n388_), .B1(new_n395_), .B2(new_n387_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n394_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n389_), .B2(KEYINPUT104), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n386_), .B1(new_n404_), .B2(new_n392_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n405_), .A2(new_n400_), .A3(new_n388_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT19), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n318_), .A2(new_n319_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n243_), .A2(new_n260_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT20), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n227_), .A2(KEYINPUT22), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT100), .B1(new_n234_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n227_), .A2(KEYINPUT22), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n229_), .A2(G169gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT100), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(G176gat), .B1(new_n415_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT101), .B1(new_n420_), .B2(new_n224_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n418_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n233_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT101), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n225_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n421_), .A2(new_n242_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n252_), .A2(new_n220_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT25), .B(G183gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n244_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n251_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n430_), .A2(new_n241_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n411_), .B1(new_n427_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n409_), .B1(new_n413_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n243_), .A2(new_n260_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n410_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n427_), .A2(new_n411_), .A3(new_n434_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n409_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT20), .A4(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(KEYINPUT102), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT102), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(new_n409_), .C1(new_n413_), .C2(new_n435_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G8gat), .B(G36gat), .Z(new_n446_));
  XNOR2_X1  g245(.A(G64gat), .B(G92gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT103), .B(KEYINPUT18), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n442_), .A2(new_n450_), .A3(new_n444_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT27), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n427_), .A2(new_n434_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n410_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(KEYINPUT20), .A3(new_n440_), .A4(new_n412_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n438_), .A2(KEYINPUT20), .A3(new_n439_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(new_n440_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n455_), .B1(new_n461_), .B2(new_n450_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n452_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n381_), .A2(new_n407_), .A3(new_n456_), .A4(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n396_), .B2(new_n401_), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT33), .B(new_n400_), .C1(new_n405_), .C2(new_n388_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT105), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n395_), .B2(new_n387_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n404_), .A2(KEYINPUT105), .A3(new_n386_), .A4(new_n392_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n400_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n451_), .A2(KEYINPUT32), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n461_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n477_));
  OAI22_X1  g276(.A1(new_n454_), .A2(new_n473_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AOI221_X4 g277(.A(KEYINPUT98), .B1(new_n354_), .B2(new_n362_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n379_), .B1(new_n378_), .B2(new_n363_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n280_), .B1(new_n464_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n280_), .A2(new_n407_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n456_), .A2(new_n463_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n484_), .A2(new_n485_), .A3(new_n381_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT73), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n488_), .A2(KEYINPUT73), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(KEYINPUT73), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n490_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G1gat), .B(G8gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT77), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499_));
  INV_X1    g298(.A(G1gat), .ZN(new_n500_));
  INV_X1    g299(.A(G8gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n497_), .A2(KEYINPUT77), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(KEYINPUT77), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n505_), .A2(new_n502_), .A3(new_n499_), .A4(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n496_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n496_), .A2(new_n510_), .A3(new_n508_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n504_), .A2(new_n507_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n492_), .A2(new_n495_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT78), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n509_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n510_), .B1(new_n496_), .B2(new_n508_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n512_), .A2(KEYINPUT78), .A3(new_n513_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT79), .A3(new_n509_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n492_), .A2(KEYINPUT15), .A3(new_n495_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT15), .B1(new_n492_), .B2(new_n495_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n508_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n518_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G169gat), .B(G197gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  NOR2_X1   g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT81), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n534_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT80), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n534_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n524_), .B2(new_n530_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n542_), .A2(KEYINPUT80), .A3(KEYINPUT81), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n536_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(new_n539_), .A3(new_n537_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT81), .B1(new_n542_), .B2(KEYINPUT80), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n535_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n487_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT66), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT67), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(KEYINPUT7), .ZN(new_n553_));
  INV_X1    g352(.A(G99gat), .ZN(new_n554_));
  INV_X1    g353(.A(G106gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n553_), .B(new_n556_), .C1(new_n551_), .C2(KEYINPUT7), .ZN(new_n557_));
  NOR2_X1   g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n558_), .B(new_n551_), .C1(new_n552_), .C2(KEYINPUT7), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT6), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(G99gat), .A3(G106gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT69), .ZN(new_n567_));
  XOR2_X1   g366(.A(G85gat), .B(G92gat), .Z(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n562_), .A2(new_n564_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n568_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT69), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(new_n573_), .A3(KEYINPUT8), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT68), .B(KEYINPUT8), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n568_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n565_), .B(KEYINPUT65), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n560_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT10), .B(G99gat), .Z(new_n581_));
  AOI22_X1  g380(.A1(KEYINPUT9), .A2(new_n568_), .B1(new_n581_), .B2(new_n555_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT64), .B(G85gat), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(G92gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT9), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n582_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n577_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n580_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G57gat), .B(G64gat), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT11), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(KEYINPUT11), .ZN(new_n594_));
  XOR2_X1   g393(.A(G71gat), .B(G78gat), .Z(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n580_), .A2(new_n598_), .A3(new_n590_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(KEYINPUT12), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n591_), .A2(new_n603_), .A3(new_n599_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT70), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n608_), .A3(new_n601_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n606_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n609_), .B(new_n610_), .C1(new_n608_), .C2(new_n600_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G120gat), .B(G148gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT72), .ZN(new_n619_));
  INV_X1    g418(.A(new_n617_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n607_), .A2(new_n611_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(KEYINPUT72), .A3(new_n617_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT13), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT37), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT76), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(KEYINPUT76), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT36), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT34), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT35), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n580_), .A2(KEYINPUT74), .A3(new_n513_), .A4(new_n590_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT8), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n572_), .B1(new_n560_), .B2(new_n565_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(new_n567_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n578_), .B1(new_n642_), .B2(new_n573_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n527_), .B1(new_n643_), .B2(new_n589_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n636_), .A2(new_n637_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n639_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n643_), .A2(new_n589_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT74), .B1(new_n647_), .B2(new_n513_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n638_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n591_), .A2(new_n527_), .B1(new_n637_), .B2(new_n636_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT74), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n591_), .B2(new_n496_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n638_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n650_), .A2(new_n652_), .A3(new_n653_), .A4(new_n639_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n633_), .B1(new_n649_), .B2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT75), .B1(new_n649_), .B2(new_n654_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n632_), .A2(KEYINPUT36), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  AOI221_X4 g458(.A(KEYINPUT75), .B1(new_n659_), .B2(new_n633_), .C1(new_n649_), .C2(new_n654_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n628_), .B(new_n629_), .C1(new_n658_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n655_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n656_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n659_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n656_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n664_), .A2(KEYINPUT76), .A3(new_n627_), .A4(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n661_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(G231gat), .A2(G233gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n598_), .B(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(new_n512_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT17), .ZN(new_n672_));
  XOR2_X1   g471(.A(G127gat), .B(G155gat), .Z(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT16), .ZN(new_n674_));
  XNOR2_X1  g473(.A(G183gat), .B(G211gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n671_), .A2(new_n672_), .A3(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(KEYINPUT17), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n671_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n667_), .A2(new_n680_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n550_), .A2(new_n626_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n407_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n500_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT38), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n624_), .A2(new_n625_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT13), .B1(new_n622_), .B2(new_n623_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n549_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n680_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n658_), .A2(new_n660_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n487_), .A2(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n690_), .A2(new_n691_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G1gat), .B1(new_n696_), .B2(new_n407_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n684_), .A2(new_n685_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n686_), .A2(new_n697_), .A3(new_n698_), .ZN(G1324gat));
  NAND3_X1  g498(.A1(new_n682_), .A2(new_n501_), .A3(new_n485_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n485_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G8gat), .B1(new_n696_), .B2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT39), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT39), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(G1325gat));
  INV_X1    g506(.A(G15gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n682_), .A2(new_n708_), .A3(new_n280_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT106), .Z(new_n710_));
  INV_X1    g509(.A(new_n280_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G15gat), .B1(new_n696_), .B2(new_n711_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n712_), .A2(KEYINPUT41), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(KEYINPUT41), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n710_), .A2(new_n713_), .A3(new_n714_), .ZN(G1326gat));
  INV_X1    g514(.A(G22gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n695_), .B2(new_n381_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT42), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n682_), .A2(new_n716_), .A3(new_n381_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1327gat));
  NOR3_X1   g519(.A1(new_n689_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n550_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G29gat), .B1(new_n723_), .B2(new_n683_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n548_), .B(new_n680_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n667_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT43), .B1(new_n487_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n667_), .B(new_n729_), .C1(new_n483_), .C2(new_n486_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n726_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n725_), .B1(new_n731_), .B2(KEYINPUT44), .ZN(new_n732_));
  INV_X1    g531(.A(new_n726_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n464_), .A2(new_n482_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n711_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n484_), .A2(new_n381_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n701_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n729_), .B1(new_n738_), .B2(new_n667_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n730_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n733_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(KEYINPUT107), .A3(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT44), .B(new_n733_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n731_), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n732_), .A2(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n683_), .A2(G29gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n724_), .B1(new_n748_), .B2(new_n749_), .ZN(G1328gat));
  NAND2_X1  g549(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(G36gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n748_), .B2(new_n485_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n722_), .A2(G36gat), .A3(new_n701_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n751_), .B(new_n754_), .C1(new_n756_), .C2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n732_), .A2(new_n743_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n746_), .A2(new_n747_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G36gat), .B1(new_n763_), .B2(new_n701_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n757_), .B(new_n758_), .Z(new_n765_));
  NAND4_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n752_), .A4(new_n753_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n760_), .A2(new_n766_), .ZN(G1329gat));
  NAND2_X1  g566(.A1(new_n280_), .A2(G43gat), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n722_), .A2(new_n711_), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n763_), .A2(new_n768_), .B1(G43gat), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n748_), .A2(new_n381_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G50gat), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n722_), .A2(G50gat), .A3(new_n481_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n772_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT111), .B(new_n775_), .C1(new_n773_), .C2(G50gat), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1331gat));
  NOR2_X1   g578(.A1(new_n626_), .A2(new_n548_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n780_), .A2(new_n691_), .A3(new_n694_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(G57gat), .A3(new_n683_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n626_), .A2(new_n487_), .A3(new_n548_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n681_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n683_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787_));
  INV_X1    g586(.A(G57gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n782_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT113), .ZN(G1332gat));
  NAND2_X1  g592(.A1(new_n781_), .A2(new_n485_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G64gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT48), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n701_), .A2(G64gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n784_), .B2(new_n797_), .ZN(G1333gat));
  NAND2_X1  g597(.A1(new_n781_), .A2(new_n280_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G71gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT49), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n711_), .A2(G71gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n784_), .B2(new_n802_), .ZN(G1334gat));
  INV_X1    g602(.A(G78gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n781_), .B2(new_n381_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT50), .Z(new_n806_));
  NAND3_X1  g605(.A1(new_n785_), .A2(new_n804_), .A3(new_n381_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1335gat));
  NOR2_X1   g607(.A1(new_n692_), .A2(new_n691_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n783_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(G85gat), .B1(new_n811_), .B2(new_n683_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n780_), .A2(new_n680_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n683_), .A2(new_n583_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT114), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n812_), .B1(new_n814_), .B2(new_n816_), .ZN(G1336gat));
  NAND3_X1  g616(.A1(new_n811_), .A2(new_n585_), .A3(new_n485_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n814_), .A2(new_n485_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n585_), .ZN(G1337gat));
  AOI21_X1  g619(.A(new_n554_), .B1(new_n814_), .B2(new_n280_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n280_), .A2(new_n581_), .ZN(new_n822_));
  OR3_X1    g621(.A1(new_n810_), .A2(KEYINPUT115), .A3(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT115), .B1(new_n810_), .B2(new_n822_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n821_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g625(.A1(new_n811_), .A2(new_n555_), .A3(new_n381_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n814_), .A2(new_n381_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(G106gat), .ZN(new_n830_));
  AOI211_X1 g629(.A(KEYINPUT52), .B(new_n555_), .C1(new_n814_), .C2(new_n381_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g632(.A1(new_n485_), .A2(new_n711_), .A3(new_n407_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT55), .B1(new_n605_), .B2(new_n606_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n607_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n605_), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n606_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n605_), .A2(KEYINPUT55), .A3(new_n606_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n837_), .A3(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n841_), .A2(KEYINPUT56), .A3(new_n617_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT56), .B1(new_n841_), .B2(new_n617_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n548_), .B(new_n621_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n523_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT79), .B1(new_n522_), .B2(new_n509_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n518_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n529_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n534_), .B1(new_n848_), .B2(new_n519_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n531_), .A2(new_n534_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n622_), .A2(new_n623_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n844_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n852_), .B2(new_n692_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n854_), .B(new_n693_), .C1(new_n844_), .C2(new_n851_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n850_), .A2(new_n621_), .A3(KEYINPUT118), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT118), .B1(new_n850_), .B2(new_n621_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n841_), .A2(new_n617_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n841_), .A2(KEYINPUT56), .A3(new_n617_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n859_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n667_), .B1(new_n864_), .B2(KEYINPUT58), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT119), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(KEYINPUT58), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n868_), .B(new_n667_), .C1(new_n864_), .C2(KEYINPUT58), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n691_), .B1(new_n856_), .B2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n626_), .A2(new_n681_), .A3(new_n549_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n481_), .B(new_n834_), .C1(new_n871_), .C2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n851_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n862_), .A2(new_n863_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n621_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n880_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n854_), .B1(new_n884_), .B2(new_n693_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n852_), .A2(KEYINPUT57), .A3(new_n692_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n869_), .A2(new_n867_), .ZN(new_n887_));
  OAI22_X1  g686(.A1(new_n842_), .A2(new_n843_), .B1(new_n858_), .B2(new_n857_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n868_), .B1(new_n890_), .B2(new_n667_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n885_), .B(new_n886_), .C1(new_n887_), .C2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n680_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n876_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n895_), .A2(KEYINPUT59), .A3(new_n481_), .A4(new_n834_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n549_), .B1(new_n879_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(G113gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n548_), .A2(new_n898_), .ZN(new_n899_));
  OAI22_X1  g698(.A1(new_n897_), .A2(new_n898_), .B1(new_n877_), .B2(new_n899_), .ZN(G1340gat));
  AOI21_X1  g699(.A(new_n626_), .B1(new_n879_), .B2(new_n896_), .ZN(new_n901_));
  INV_X1    g700(.A(G120gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n626_), .B2(KEYINPUT60), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(KEYINPUT60), .B2(new_n902_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n901_), .A2(new_n902_), .B1(new_n877_), .B2(new_n904_), .ZN(G1341gat));
  INV_X1    g704(.A(G127gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n877_), .B2(new_n680_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT120), .B(new_n906_), .C1(new_n877_), .C2(new_n680_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n879_), .A2(new_n896_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n691_), .A2(G127gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT121), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n909_), .A2(new_n910_), .B1(new_n911_), .B2(new_n913_), .ZN(G1342gat));
  INV_X1    g713(.A(G134gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n877_), .B2(new_n692_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  OAI211_X1 g717(.A(KEYINPUT122), .B(new_n915_), .C1(new_n877_), .C2(new_n692_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT123), .B(G134gat), .Z(new_n920_));
  NOR2_X1   g719(.A1(new_n727_), .A2(new_n920_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n918_), .A2(new_n919_), .B1(new_n911_), .B2(new_n921_), .ZN(G1343gat));
  AOI21_X1  g721(.A(new_n876_), .B1(new_n892_), .B2(new_n680_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n280_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n485_), .A2(new_n481_), .A3(new_n407_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  OR3_X1    g725(.A1(new_n926_), .A2(G141gat), .A3(new_n549_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G141gat), .B1(new_n926_), .B2(new_n549_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1344gat));
  OR3_X1    g728(.A1(new_n926_), .A2(G148gat), .A3(new_n626_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G148gat), .B1(new_n926_), .B2(new_n626_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1345gat));
  XNOR2_X1  g731(.A(KEYINPUT61), .B(G155gat), .ZN(new_n933_));
  OR3_X1    g732(.A1(new_n926_), .A2(new_n680_), .A3(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n926_), .B2(new_n680_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1346gat));
  OAI21_X1  g735(.A(G162gat), .B1(new_n926_), .B2(new_n727_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n693_), .A2(new_n332_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n926_), .B2(new_n938_), .ZN(G1347gat));
  NOR2_X1   g738(.A1(new_n701_), .A2(new_n484_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n549_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n481_), .B(new_n942_), .C1(new_n871_), .C2(new_n876_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(G169gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(KEYINPUT125), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n943_), .A2(new_n946_), .A3(G169gat), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n945_), .A2(new_n947_), .A3(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n422_), .A2(new_n423_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n943_), .A2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n946_), .B1(new_n943_), .B2(G169gat), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(new_n948_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n950_), .A2(new_n954_), .ZN(G1348gat));
  NAND3_X1  g754(.A1(new_n895_), .A2(new_n481_), .A3(new_n940_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(G176gat), .B1(new_n957_), .B2(new_n689_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n956_), .A2(new_n233_), .A3(new_n626_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1349gat));
  NOR3_X1   g759(.A1(new_n956_), .A2(new_n431_), .A3(new_n680_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n957_), .A2(new_n691_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n961_), .B1(new_n245_), .B2(new_n962_), .ZN(G1350gat));
  OAI21_X1  g762(.A(G190gat), .B1(new_n956_), .B2(new_n727_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n693_), .A2(new_n244_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n964_), .B1(new_n956_), .B2(new_n965_), .ZN(G1351gat));
  NOR3_X1   g765(.A1(new_n701_), .A2(new_n481_), .A3(new_n683_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n924_), .A2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n309_), .B1(new_n968_), .B2(new_n549_), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n924_), .A2(G197gat), .A3(new_n548_), .A4(new_n967_), .ZN(new_n970_));
  AND2_X1   g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1352gat));
  AND2_X1   g770(.A1(new_n924_), .A2(new_n967_), .ZN(new_n972_));
  OAI211_X1 g771(.A(new_n972_), .B(new_n689_), .C1(KEYINPUT126), .C2(new_n310_), .ZN(new_n973_));
  XOR2_X1   g772(.A(KEYINPUT126), .B(G204gat), .Z(new_n974_));
  OAI21_X1  g773(.A(new_n974_), .B1(new_n968_), .B2(new_n626_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n975_), .ZN(G1353gat));
  XNOR2_X1  g775(.A(KEYINPUT63), .B(G211gat), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n972_), .A2(new_n691_), .A3(new_n977_), .ZN(new_n978_));
  OAI22_X1  g777(.A1(new_n968_), .A2(new_n680_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n978_), .A2(new_n979_), .ZN(G1354gat));
  NAND2_X1  g779(.A1(new_n667_), .A2(G218gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(KEYINPUT127), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n924_), .A2(new_n693_), .A3(new_n967_), .ZN(new_n983_));
  INV_X1    g782(.A(G218gat), .ZN(new_n984_));
  AOI22_X1  g783(.A1(new_n972_), .A2(new_n982_), .B1(new_n983_), .B2(new_n984_), .ZN(G1355gat));
endmodule


