//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203_));
  INV_X1    g002(.A(G36gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G29gat), .ZN(new_n205_));
  INV_X1    g004(.A(G29gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G36gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT71), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT71), .B1(new_n205_), .B2(new_n207_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT72), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT71), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n206_), .A2(G36gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n204_), .A2(G29gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT72), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT71), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n210_), .A2(new_n211_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n211_), .B1(new_n210_), .B2(new_n218_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n203_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n225_), .A3(KEYINPUT65), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT9), .ZN(new_n232_));
  AND2_X1   g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G85gat), .A2(G92gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n232_), .B1(new_n235_), .B2(KEYINPUT9), .ZN(new_n236_));
  OR2_X1    g035(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n240_), .A2(new_n241_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n230_), .B(new_n236_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n245_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n246_));
  INV_X1    g045(.A(G85gat), .ZN(new_n247_));
  INV_X1    g046(.A(G92gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT67), .A3(new_n231_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT8), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G99gat), .A2(G106gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT7), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT66), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n259_), .A3(new_n256_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n254_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n252_), .B1(new_n230_), .B2(new_n261_), .ZN(new_n262_));
  NOR4_X1   g061(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n259_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n226_), .B(new_n253_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n246_), .A2(new_n250_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n251_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n244_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n211_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT72), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n216_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n210_), .A2(new_n218_), .A3(new_n211_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(KEYINPUT15), .A3(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n221_), .A2(new_n268_), .A3(new_n274_), .ZN(new_n275_));
  OAI221_X1 g074(.A(new_n244_), .B1(new_n262_), .B2(new_n267_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G232gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT34), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT35), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .A4(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n281_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n275_), .A2(new_n284_), .A3(new_n276_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n282_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n275_), .B2(KEYINPUT73), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n283_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G190gat), .B(G218gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G134gat), .B(G162gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT36), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(KEYINPUT36), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n288_), .B2(new_n295_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n293_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT37), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT76), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(KEYINPUT76), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n288_), .A2(new_n295_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n294_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n307_), .A2(KEYINPUT76), .A3(new_n299_), .A4(new_n293_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G15gat), .B(G22gat), .ZN(new_n310_));
  INV_X1    g109(.A(G1gat), .ZN(new_n311_));
  INV_X1    g110(.A(G8gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT14), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G8gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G64gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G57gat), .ZN(new_n320_));
  INV_X1    g119(.A(G57gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G64gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT11), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G71gat), .B(G78gat), .Z(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n323_), .A2(KEYINPUT68), .A3(new_n324_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT68), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G57gat), .B(G64gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(KEYINPUT11), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n327_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT68), .B1(new_n323_), .B2(new_n324_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n329_), .A3(KEYINPUT11), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(new_n325_), .A3(new_n334_), .A4(new_n326_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n318_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT17), .ZN(new_n338_));
  XOR2_X1   g137(.A(G127gat), .B(G155gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G183gat), .B(G211gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n337_), .A2(new_n338_), .A3(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(KEYINPUT17), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n337_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n309_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G120gat), .B(G148gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT5), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G176gat), .B(G204gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT70), .ZN(new_n353_));
  INV_X1    g152(.A(new_n336_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n268_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n336_), .B(new_n244_), .C1(new_n262_), .C2(new_n267_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G230gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(KEYINPUT69), .A3(new_n359_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n355_), .A2(KEYINPUT12), .A3(new_n356_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT12), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n268_), .A2(new_n354_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n359_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n353_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n367_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n358_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n371_), .A2(new_n362_), .A3(new_n363_), .A4(new_n352_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT13), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n348_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT78), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n377_));
  AOI21_X1  g176(.A(G176gat), .B1(new_n377_), .B2(KEYINPUT22), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G169gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n381_), .A2(KEYINPUT23), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n379_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT25), .B(G183gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT24), .A3(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n391_), .A2(KEYINPUT24), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n380_), .A2(KEYINPUT23), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n383_), .B2(new_n380_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n387_), .A2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n399_), .B(KEYINPUT30), .Z(new_n400_));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(G15gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G71gat), .ZN(new_n404_));
  INV_X1    g203(.A(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n400_), .B(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G127gat), .B(G134gat), .Z(new_n409_));
  XOR2_X1   g208(.A(G113gat), .B(G120gat), .Z(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n408_), .A2(new_n412_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(G43gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT31), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT84), .ZN(new_n424_));
  NOR3_X1   g223(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT86), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G141gat), .A2(G148gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT87), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT2), .ZN(new_n429_));
  OR2_X1    g228(.A1(G141gat), .A2(G148gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT3), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT2), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n427_), .A2(KEYINPUT87), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n424_), .B1(new_n426_), .B2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n430_), .A2(new_n427_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT1), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G155gat), .A2(G162gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n441_));
  OR3_X1    g240(.A1(new_n439_), .A2(new_n441_), .A3(KEYINPUT1), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n439_), .B2(KEYINPUT1), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n424_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n436_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n445_), .A3(new_n412_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n439_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n445_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n411_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(KEYINPUT4), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G225gat), .A2(G233gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT96), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n440_), .A2(new_n445_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n411_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n451_), .A2(new_n454_), .A3(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G29gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G85gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT0), .B(G57gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n446_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n384_), .A2(new_n393_), .A3(new_n394_), .A4(new_n390_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n392_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G169gat), .ZN(new_n469_));
  INV_X1    g268(.A(G176gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT93), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n397_), .B2(new_n386_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n471_), .A2(KEYINPUT93), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n467_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G197gat), .A2(G204gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT88), .B(G204gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(G197gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT89), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G211gat), .B(G218gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT21), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n478_), .A2(KEYINPUT89), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n478_), .A2(KEYINPUT21), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n477_), .A2(G197gat), .ZN(new_n486_));
  INV_X1    g285(.A(G197gat), .ZN(new_n487_));
  INV_X1    g286(.A(G204gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT21), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n480_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  OAI22_X1  g289(.A1(new_n483_), .A2(new_n484_), .B1(new_n485_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n466_), .B1(new_n475_), .B2(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n478_), .A2(KEYINPUT89), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n494_));
  OAI221_X1 g293(.A(new_n480_), .B1(new_n486_), .B2(new_n489_), .C1(KEYINPUT21), .C2(new_n478_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n387_), .A3(new_n495_), .A4(new_n398_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G226gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT19), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G8gat), .B(G36gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G64gat), .B(G92gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n399_), .A2(new_n491_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n474_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n397_), .A2(new_n386_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n472_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n509_), .A2(new_n494_), .A3(new_n495_), .A4(new_n467_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n499_), .A2(new_n466_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n506_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n500_), .A2(new_n505_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n505_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n499_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n506_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n514_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n513_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n465_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n451_), .A2(new_n453_), .A3(new_n457_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n446_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n462_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(KEYINPUT33), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n525_), .B(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT98), .B1(new_n522_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n527_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n525_), .B(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n505_), .B1(new_n500_), .B2(new_n512_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n516_), .A2(new_n517_), .A3(new_n514_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT95), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n513_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT98), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n531_), .A2(new_n536_), .A3(new_n537_), .A4(new_n465_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n523_), .A2(new_n524_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n463_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(KEYINPUT100), .A3(new_n525_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT100), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n539_), .A2(new_n542_), .A3(new_n463_), .ZN(new_n543_));
  OR2_X1    g342(.A1(KEYINPUT99), .A2(KEYINPUT20), .ZN(new_n544_));
  NAND2_X1  g343(.A1(KEYINPUT99), .A2(KEYINPUT20), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n510_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n506_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n499_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n499_), .B2(new_n497_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT32), .A3(new_n505_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n505_), .A2(KEYINPUT32), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n500_), .A2(new_n512_), .A3(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n541_), .A2(new_n543_), .A3(new_n550_), .A4(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n529_), .A2(new_n538_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G228gat), .A2(G233gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT29), .B1(new_n448_), .B2(new_n449_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n491_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n556_), .A3(new_n491_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G78gat), .B(G106gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n559_), .A2(KEYINPUT91), .A3(new_n560_), .A4(new_n562_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n560_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n561_), .B1(new_n568_), .B2(new_n558_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT28), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n448_), .A2(new_n449_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT29), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR4_X1   g373(.A1(new_n448_), .A2(new_n449_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G22gat), .B(G50gat), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n577_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n567_), .A2(new_n569_), .A3(new_n578_), .A4(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n555_), .B1(new_n566_), .B2(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n569_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n583_), .A2(KEYINPUT92), .A3(new_n565_), .A4(new_n567_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT90), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n569_), .A2(new_n563_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n578_), .A2(new_n580_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n587_), .B(new_n588_), .C1(new_n586_), .C2(new_n569_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n554_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n541_), .A2(new_n543_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n549_), .A2(new_n514_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(KEYINPUT27), .A3(new_n513_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT27), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n422_), .B1(new_n591_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n422_), .A2(new_n592_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n585_), .A2(new_n589_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n599_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n316_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT79), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n272_), .A2(new_n273_), .A3(new_n316_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n272_), .A2(KEYINPUT79), .A3(new_n273_), .A4(new_n316_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n221_), .A2(new_n274_), .A3(new_n316_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n612_), .A3(new_n608_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT80), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G169gat), .B(G197gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n618_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n615_), .A2(new_n617_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n376_), .A2(new_n606_), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n311_), .A3(new_n593_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n606_), .A2(new_n298_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n374_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n631_), .A2(new_n347_), .A3(new_n627_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n592_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n202_), .B1(new_n629_), .B2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n202_), .B2(new_n629_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1324gat));
  NAND3_X1  g437(.A1(new_n628_), .A2(new_n312_), .A3(new_n599_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n633_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n599_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642_));
  AND4_X1   g441(.A1(KEYINPUT102), .A2(new_n641_), .A3(new_n642_), .A4(G8gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n312_), .B1(new_n644_), .B2(KEYINPUT39), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n641_), .A2(new_n645_), .B1(KEYINPUT102), .B2(new_n642_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n639_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n639_), .B(new_n648_), .C1(new_n643_), .C2(new_n646_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1325gat));
  AOI21_X1  g451(.A(new_n402_), .B1(new_n640_), .B2(new_n422_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT41), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n628_), .A2(new_n402_), .A3(new_n422_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1326gat));
  OAI21_X1  g455(.A(G22gat), .B1(new_n633_), .B2(new_n590_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n628_), .A2(new_n659_), .A3(new_n604_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(new_n298_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n347_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n374_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n626_), .B(new_n666_), .C1(new_n602_), .C2(new_n605_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT107), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n604_), .A2(new_n599_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n592_), .A3(new_n422_), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n554_), .A2(new_n590_), .B1(new_n594_), .B2(new_n600_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n422_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n626_), .A4(new_n666_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n668_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n593_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n374_), .A2(new_n347_), .A3(new_n626_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT104), .Z(new_n679_));
  NAND2_X1  g478(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n309_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n606_), .B2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n309_), .B(new_n680_), .C1(new_n602_), .C2(new_n605_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n679_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n677_), .B1(new_n688_), .B2(KEYINPUT44), .ZN(new_n689_));
  INV_X1    g488(.A(new_n679_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n687_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n683_), .B1(new_n672_), .B2(new_n309_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(KEYINPUT106), .A3(new_n694_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n689_), .A2(new_n695_), .B1(KEYINPUT44), .B2(new_n688_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n592_), .A2(new_n206_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n676_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(KEYINPUT108), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n688_), .A2(KEYINPUT44), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n688_), .A2(new_n677_), .A3(KEYINPUT44), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT106), .B1(new_n693_), .B2(new_n694_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n599_), .B(new_n702_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n600_), .A2(G36gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n668_), .A2(new_n674_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT45), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n668_), .A2(new_n710_), .A3(new_n674_), .A4(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n699_), .A2(KEYINPUT108), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n701_), .B1(new_n706_), .B2(new_n715_), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n700_), .B(new_n714_), .C1(new_n705_), .C2(G36gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  AOI21_X1  g517(.A(G43gat), .B1(new_n675_), .B2(new_n422_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n422_), .A2(G43gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n696_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n675_), .B2(new_n604_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n604_), .A2(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n696_), .B2(new_n725_), .ZN(G1331gat));
  NOR3_X1   g525(.A1(new_n374_), .A2(new_n347_), .A3(new_n626_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n630_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n592_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n374_), .A2(new_n626_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n672_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n348_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n593_), .A2(new_n321_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(G1332gat));
  OAI21_X1  g533(.A(G64gat), .B1(new_n728_), .B2(new_n600_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n732_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n319_), .A3(new_n599_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741_));
  INV_X1    g540(.A(new_n728_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n422_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n738_), .A2(new_n741_), .A3(new_n422_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1334gat));
  OAI21_X1  g546(.A(G78gat), .B1(new_n728_), .B2(new_n590_), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n590_), .A2(G78gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n732_), .B2(new_n751_), .ZN(G1335gat));
  NAND2_X1  g551(.A1(new_n731_), .A2(new_n664_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n247_), .A3(new_n593_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n730_), .A2(new_n347_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT112), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n593_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n760_), .B2(new_n247_), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n754_), .A2(new_n248_), .A3(new_n599_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n759_), .A2(new_n599_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n248_), .ZN(G1337gat));
  NAND4_X1  g563(.A1(new_n754_), .A2(new_n422_), .A3(new_n237_), .A4(new_n239_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n759_), .A2(new_n422_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n405_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(KEYINPUT113), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n767_), .B(new_n769_), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n754_), .A2(new_n238_), .A3(new_n604_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n759_), .A2(new_n604_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(G106gat), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT52), .B(new_n238_), .C1(new_n759_), .C2(new_n604_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g576(.A(new_n592_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n669_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(KEYINPUT59), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT54), .B1(new_n375_), .B2(new_n626_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n348_), .A2(new_n783_), .A3(new_n627_), .A4(new_n374_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n626_), .A2(new_n372_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n358_), .A2(KEYINPUT114), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(new_n788_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n371_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n370_), .A2(KEYINPUT55), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n353_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n787_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n789_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n368_), .B2(new_n791_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n353_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n786_), .B1(new_n796_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n616_), .A2(new_n608_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n616_), .A2(KEYINPUT115), .A3(new_n608_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n613_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n611_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n622_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n625_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n802_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n662_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n662_), .B(KEYINPUT57), .C1(new_n802_), .C2(new_n812_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n372_), .A3(new_n625_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n796_), .B2(new_n801_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(KEYINPUT116), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n823_), .B(new_n820_), .C1(new_n796_), .C2(new_n801_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n309_), .B(new_n818_), .C1(new_n822_), .C2(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n810_), .A2(new_n372_), .A3(new_n625_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n793_), .A2(new_n795_), .A3(new_n787_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n800_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n829_), .A2(KEYINPUT118), .A3(new_n819_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n821_), .B2(KEYINPUT58), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n825_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n823_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n821_), .A2(KEYINPUT116), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n819_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n818_), .B1(new_n837_), .B2(new_n309_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n817_), .B1(new_n834_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n347_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n785_), .B1(KEYINPUT121), .B2(new_n840_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n840_), .A2(KEYINPUT121), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n781_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT122), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(G113gat), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n844_), .A2(G113gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n626_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n839_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n817_), .B(KEYINPUT119), .C1(new_n834_), .C2(new_n838_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n347_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n785_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n779_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT120), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n663_), .B1(new_n839_), .B2(new_n848_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n785_), .B1(new_n857_), .B2(new_n850_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n856_), .B(KEYINPUT59), .C1(new_n858_), .C2(new_n779_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n843_), .B(new_n847_), .C1(new_n855_), .C2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G113gat), .B1(new_n853_), .B2(new_n626_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT123), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n855_), .A2(new_n859_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n843_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n847_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  INV_X1    g666(.A(new_n861_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n862_), .A2(new_n869_), .ZN(G1340gat));
  AOI21_X1  g669(.A(new_n843_), .B1(new_n855_), .B2(new_n859_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n871_), .A2(new_n631_), .ZN(new_n872_));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n853_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n374_), .B2(KEYINPUT60), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(KEYINPUT60), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(KEYINPUT124), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(KEYINPUT124), .B2(new_n875_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n872_), .A2(new_n873_), .B1(new_n874_), .B2(new_n878_), .ZN(G1341gat));
  AOI21_X1  g678(.A(G127gat), .B1(new_n853_), .B2(new_n663_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT125), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n663_), .A2(G127gat), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT126), .Z(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n871_), .B2(new_n883_), .ZN(G1342gat));
  INV_X1    g683(.A(G134gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n853_), .A2(new_n885_), .A3(new_n298_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n871_), .A2(new_n309_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1343gat));
  INV_X1    g687(.A(new_n858_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n422_), .A2(new_n599_), .A3(new_n592_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n604_), .A3(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n627_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n374_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT127), .B(G148gat), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1345gat));
  NOR2_X1   g695(.A1(new_n891_), .A2(new_n347_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT61), .B(G155gat), .Z(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n891_), .B2(new_n685_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n662_), .A2(G162gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n891_), .B2(new_n901_), .ZN(G1347gat));
  AOI21_X1  g701(.A(new_n604_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n603_), .A2(new_n600_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905_), .B2(new_n627_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n905_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n469_), .A3(new_n626_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT62), .B(G169gat), .C1(new_n905_), .C2(new_n627_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n908_), .A2(new_n910_), .A3(new_n911_), .ZN(G1348gat));
  AOI21_X1  g711(.A(G176gat), .B1(new_n909_), .B2(new_n631_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n858_), .A2(new_n604_), .ZN(new_n914_));
  NOR4_X1   g713(.A1(new_n603_), .A2(new_n470_), .A3(new_n600_), .A4(new_n374_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n663_), .A3(new_n904_), .ZN(new_n917_));
  INV_X1    g716(.A(G183gat), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n603_), .A2(new_n388_), .A3(new_n600_), .A4(new_n347_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n917_), .A2(new_n918_), .B1(new_n903_), .B2(new_n919_), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n905_), .B2(new_n685_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n298_), .A2(new_n389_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n905_), .B2(new_n922_), .ZN(G1351gat));
  NOR4_X1   g722(.A1(new_n590_), .A2(new_n422_), .A3(new_n593_), .A4(new_n600_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n889_), .A2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n627_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n487_), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n374_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(G204gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n477_), .B2(new_n928_), .ZN(G1353gat));
  INV_X1    g729(.A(new_n925_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n663_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AND2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n932_), .B2(new_n933_), .ZN(G1354gat));
  OR3_X1    g735(.A1(new_n925_), .A2(G218gat), .A3(new_n662_), .ZN(new_n937_));
  OAI21_X1  g736(.A(G218gat), .B1(new_n925_), .B2(new_n685_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1355gat));
endmodule


