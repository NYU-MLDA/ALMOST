//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT9), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n208_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  OR3_X1    g022(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n217_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n206_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT65), .B1(new_n227_), .B2(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  AOI211_X1 g029(.A(new_n229_), .B(new_n230_), .C1(new_n226_), .C2(new_n206_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n209_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n230_), .A3(new_n206_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n214_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT15), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G29gat), .B(G36gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G43gat), .B(G50gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n236_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT15), .A3(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n235_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n242_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(new_n235_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G232gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT34), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n245_), .A2(new_n247_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n227_), .A2(KEYINPUT8), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n229_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n227_), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n234_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n213_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n251_), .A2(KEYINPUT35), .A3(new_n253_), .A4(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n253_), .A2(KEYINPUT35), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT35), .B(new_n253_), .C1(new_n249_), .C2(KEYINPUT71), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n243_), .A2(new_n244_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n260_), .B1(new_n266_), .B2(new_n259_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G190gat), .B(G218gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G134gat), .ZN(new_n271_));
  INV_X1    g070(.A(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT36), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n202_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n269_), .A2(new_n202_), .A3(new_n275_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n273_), .B(KEYINPUT36), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n263_), .A2(new_n264_), .A3(new_n268_), .A4(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT37), .B1(new_n279_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n278_), .ZN(new_n287_));
  OAI211_X1 g086(.A(KEYINPUT37), .B(new_n281_), .C1(new_n287_), .C2(new_n276_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT74), .B(G1gat), .Z(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G8gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n295_), .B(G1gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G57gat), .B(G64gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n302_), .A2(KEYINPUT11), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(KEYINPUT11), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G71gat), .B(G78gat), .ZN(new_n305_));
  OR3_X1    g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n305_), .A3(KEYINPUT11), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G231gat), .A2(G233gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT75), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n308_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n301_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT17), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT16), .B(G183gat), .ZN(new_n315_));
  INV_X1    g114(.A(G211gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G155gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n313_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n314_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n312_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n290_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT76), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT19), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G169gat), .ZN(new_n330_));
  INV_X1    g129(.A(G176gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n332_), .A2(KEYINPUT84), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT23), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT83), .B(G190gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(G183gat), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(KEYINPUT84), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G169gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n331_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT24), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT24), .A3(new_n328_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n335_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n336_), .A2(KEYINPUT26), .ZN(new_n345_));
  NOR2_X1   g144(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT81), .B(KEYINPUT25), .ZN(new_n351_));
  INV_X1    g150(.A(G183gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(KEYINPUT82), .B(new_n350_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT82), .B1(new_n351_), .B2(G183gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n344_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n339_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G197gat), .B(G204gat), .Z(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT21), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G197gat), .B(G204gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT21), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT90), .ZN(new_n363_));
  INV_X1    g162(.A(G218gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n316_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G211gat), .A2(G218gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n363_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n359_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(KEYINPUT21), .A3(new_n358_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT20), .B1(new_n357_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  OR2_X1    g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n335_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n332_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT94), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n379_));
  NAND2_X1  g178(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n340_), .A3(new_n331_), .ZN(new_n382_));
  AND2_X1   g181(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n383_));
  AND2_X1   g182(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n384_));
  OAI22_X1  g183(.A1(new_n349_), .A2(new_n383_), .B1(new_n384_), .B2(new_n346_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n379_), .A2(new_n341_), .A3(new_n380_), .A4(new_n328_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT93), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT93), .B1(new_n385_), .B2(new_n386_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n382_), .B(new_n335_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n373_), .B1(new_n378_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n327_), .B1(new_n372_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n378_), .A2(new_n373_), .A3(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n357_), .A2(new_n371_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n327_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(KEYINPUT20), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT18), .B(G64gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G92gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  XNOR2_X1  g199(.A(new_n396_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n368_), .A2(KEYINPUT91), .A3(new_n370_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT91), .B1(new_n368_), .B2(new_n370_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n389_), .B(new_n376_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n393_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT98), .B1(new_n407_), .B2(KEYINPUT20), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n327_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n372_), .A2(new_n390_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n394_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n412_), .B(new_n327_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n400_), .B(KEYINPUT101), .Z(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT102), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n391_), .A2(new_n400_), .A3(new_n395_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n415_), .A2(KEYINPUT102), .A3(new_n416_), .A4(new_n417_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n404_), .B1(new_n423_), .B2(KEYINPUT27), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G127gat), .B(G134gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G113gat), .B(G120gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n427_), .A2(new_n429_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n436_), .B(KEYINPUT3), .Z(new_n437_));
  NAND2_X1  g236(.A1(G141gat), .A2(G148gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n438_), .B(KEYINPUT2), .Z(new_n439_));
  OAI21_X1  g238(.A(new_n435_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n436_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(KEYINPUT1), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n438_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n432_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n447_), .A2(KEYINPUT4), .A3(new_n448_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n430_), .A2(new_n431_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(KEYINPUT95), .A3(new_n455_), .A4(new_n445_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n451_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n448_), .B2(KEYINPUT4), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n453_), .A2(new_n456_), .A3(new_n457_), .A4(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n452_), .A2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G1gat), .B(G29gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT97), .ZN(new_n463_));
  XOR2_X1   g262(.A(G57gat), .B(G85gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n461_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(new_n452_), .A3(new_n460_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(KEYINPUT100), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT100), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n461_), .A2(new_n472_), .A3(new_n467_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n445_), .A2(KEYINPUT29), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n475_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G228gat), .A2(G233gat), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(KEYINPUT89), .Z(new_n479_));
  OR3_X1    g278(.A1(new_n475_), .A2(new_n373_), .A3(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G22gat), .B(G50gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G78gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n480_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n445_), .A2(KEYINPUT29), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT28), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(new_n204_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n489_), .B(G106gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n357_), .A2(KEYINPUT30), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT30), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n339_), .A2(new_n356_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G15gat), .B(G43gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n495_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT85), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  NAND3_X1  g305(.A1(new_n500_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT88), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n507_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n432_), .B(KEYINPUT31), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(KEYINPUT88), .B(new_n514_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n474_), .A2(new_n494_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT103), .B1(new_n424_), .B2(new_n518_), .ZN(new_n519_));
  AND4_X1   g318(.A1(new_n474_), .A2(new_n494_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT103), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n422_), .A2(new_n421_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n402_), .B1(new_n522_), .B2(new_n420_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n520_), .B(new_n521_), .C1(new_n523_), .C2(new_n404_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n423_), .A2(KEYINPUT27), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n494_), .B1(new_n525_), .B2(new_n403_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n470_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(KEYINPUT33), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n450_), .A2(new_n457_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n453_), .A2(new_n459_), .A3(new_n456_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n529_), .B(new_n467_), .C1(new_n530_), .C2(new_n457_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(KEYINPUT33), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n528_), .A2(new_n531_), .A3(new_n401_), .A4(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n415_), .A2(KEYINPUT32), .A3(new_n400_), .A4(new_n416_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n400_), .A2(KEYINPUT32), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n391_), .A2(new_n535_), .A3(new_n395_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n471_), .A2(new_n534_), .A3(new_n473_), .A4(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n526_), .A2(new_n474_), .B1(new_n538_), .B2(new_n494_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n516_), .A2(new_n517_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n519_), .B(new_n524_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n235_), .B2(new_n308_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n235_), .B2(new_n308_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n308_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n259_), .A2(KEYINPUT12), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n543_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT67), .B(G204gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G120gat), .B(G148gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT5), .B(G176gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT66), .B1(new_n259_), .B2(new_n547_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT66), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n235_), .A2(new_n556_), .A3(new_n308_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n259_), .A2(new_n547_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n549_), .B(new_n554_), .C1(new_n560_), .C2(new_n544_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n554_), .B(KEYINPUT68), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n544_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n549_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT13), .Z(new_n567_));
  NAND3_X1  g366(.A1(new_n254_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n266_), .A2(KEYINPUT77), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT77), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n250_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n301_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT78), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT79), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n572_), .A2(new_n301_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n569_), .A2(new_n571_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n580_));
  OAI211_X1 g379(.A(G229gat), .B(G233gat), .C1(new_n579_), .C2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n568_), .A2(new_n573_), .A3(KEYINPUT79), .A4(new_n575_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n340_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(G197gat), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(KEYINPUT80), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n583_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n567_), .A2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n541_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n325_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n474_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n291_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT38), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n277_), .A2(new_n278_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n591_), .A2(new_n323_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(KEYINPUT104), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n600_), .B(new_n541_), .C1(KEYINPUT104), .C2(new_n599_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n474_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(G1324gat));
  INV_X1    g402(.A(new_n424_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G8gat), .B1(new_n601_), .B2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(KEYINPUT105), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT39), .B1(new_n605_), .B2(KEYINPUT105), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  NAND3_X1  g407(.A1(new_n594_), .A2(new_n292_), .A3(new_n424_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(G1325gat));
  INV_X1    g411(.A(new_n540_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G15gat), .B1(new_n601_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT41), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n593_), .A2(G15gat), .A3(new_n613_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1326gat));
  OAI21_X1  g416(.A(G22gat), .B1(new_n601_), .B2(new_n494_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT42), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n494_), .A2(G22gat), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n593_), .B2(new_n620_), .ZN(G1327gat));
  INV_X1    g420(.A(new_n323_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n598_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT107), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n592_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(G29gat), .B1(new_n626_), .B2(new_n595_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n288_), .B1(new_n598_), .B2(KEYINPUT37), .ZN(new_n628_));
  INV_X1    g427(.A(new_n494_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n474_), .B(new_n629_), .C1(new_n523_), .C2(new_n404_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n538_), .A2(new_n494_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n540_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n519_), .A2(new_n524_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n628_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n628_), .B2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n634_), .A2(new_n637_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n591_), .B(new_n622_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n634_), .B(new_n637_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(KEYINPUT44), .A3(new_n591_), .A4(new_n622_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(G29gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n627_), .B1(new_n646_), .B2(new_n595_), .ZN(G1328gat));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT109), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n642_), .A2(new_n644_), .A3(new_n424_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT108), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT108), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n653_), .A3(G36gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n625_), .A2(G36gat), .A3(new_n604_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT45), .Z(new_n657_));
  AOI21_X1  g456(.A(new_n649_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n650_), .A2(new_n653_), .A3(G36gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n653_), .B1(new_n650_), .B2(G36gat), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n657_), .B(new_n649_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n648_), .B1(new_n658_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT109), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(KEYINPUT46), .A3(new_n661_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(G1329gat));
  NAND3_X1  g466(.A1(new_n645_), .A2(G43gat), .A3(new_n540_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT110), .B(G43gat), .Z(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n625_), .B2(new_n613_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g471(.A(G50gat), .B1(new_n626_), .B2(new_n629_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n629_), .A2(G50gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n645_), .B2(new_n674_), .ZN(G1331gat));
  INV_X1    g474(.A(new_n567_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n589_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n541_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n325_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G57gat), .B1(new_n680_), .B2(new_n595_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n323_), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n598_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n681_), .B1(new_n684_), .B2(new_n595_), .ZN(G1332gat));
  OR3_X1    g484(.A1(new_n679_), .A2(G64gat), .A3(new_n604_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n682_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n598_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n424_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G64gat), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT48), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT48), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n686_), .B1(new_n691_), .B2(new_n692_), .ZN(G1333gat));
  OR3_X1    g492(.A1(new_n679_), .A2(G71gat), .A3(new_n613_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n687_), .A2(new_n688_), .A3(new_n540_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G71gat), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT49), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT49), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1334gat));
  OR3_X1    g498(.A1(new_n679_), .A2(G78gat), .A3(new_n494_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n687_), .A2(new_n688_), .A3(new_n629_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G78gat), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT50), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT50), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1335gat));
  NAND2_X1  g504(.A1(new_n678_), .A2(new_n624_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n210_), .B1(new_n706_), .B2(new_n474_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT111), .Z(new_n708_));
  AND3_X1   g507(.A1(new_n643_), .A2(new_n622_), .A3(new_n677_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n474_), .A2(new_n210_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n709_), .B2(new_n710_), .ZN(G1336gat));
  NAND3_X1  g510(.A1(new_n709_), .A2(G92gat), .A3(new_n424_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n211_), .B1(new_n706_), .B2(new_n604_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1337gat));
  INV_X1    g513(.A(new_n203_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n706_), .A2(new_n715_), .A3(new_n613_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n709_), .A2(new_n540_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(G99gat), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g518(.A(new_n204_), .B1(new_n709_), .B2(new_n629_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT52), .Z(new_n721_));
  NOR3_X1   g520(.A1(new_n706_), .A2(G106gat), .A3(new_n494_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT112), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g524(.A(G113gat), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n613_), .A2(new_n474_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n604_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n549_), .A2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n543_), .A2(new_n546_), .A3(KEYINPUT55), .A4(new_n548_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n543_), .A2(new_n548_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n544_), .B1(new_n734_), .B2(new_n558_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n562_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n556_), .B1(new_n235_), .B2(new_n308_), .ZN(new_n739_));
  AND4_X1   g538(.A1(new_n556_), .A2(new_n258_), .A3(new_n213_), .A4(new_n308_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n543_), .A2(new_n548_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n545_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n562_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n738_), .A2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n578_), .A2(new_n587_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n575_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n579_), .A2(new_n580_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n575_), .B1(new_n568_), .B2(new_n573_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n586_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n747_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n561_), .A3(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(KEYINPUT58), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n753_), .B(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n756_), .A2(new_n290_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n738_), .A2(new_n758_), .A3(new_n745_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n561_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n562_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(KEYINPUT113), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(new_n589_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n759_), .A2(new_n762_), .A3(KEYINPUT114), .A4(new_n589_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n752_), .A2(new_n566_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n765_), .A2(new_n766_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n688_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(new_n688_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n757_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n770_), .A2(new_n688_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n775_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n770_), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n688_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n323_), .B1(new_n776_), .B2(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n290_), .A2(new_n590_), .A3(new_n676_), .A4(new_n323_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT54), .Z(new_n784_));
  OAI211_X1 g583(.A(new_n494_), .B(new_n729_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT59), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(KEYINPUT120), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(KEYINPUT120), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n778_), .A2(KEYINPUT116), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n770_), .A2(new_n771_), .A3(new_n688_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n775_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n757_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n779_), .A4(new_n780_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n622_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n784_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n629_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n792_), .B1(new_n800_), .B2(new_n729_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n726_), .B1(new_n790_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n800_), .B2(new_n729_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n784_), .B1(new_n797_), .B2(new_n622_), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n806_), .A2(KEYINPUT119), .A3(new_n629_), .A4(new_n728_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n589_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n803_), .A2(new_n589_), .B1(new_n726_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n676_), .B2(KEYINPUT60), .ZN(new_n811_));
  OAI221_X1 g610(.A(new_n811_), .B1(KEYINPUT60), .B2(new_n810_), .C1(new_n805_), .C2(new_n807_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n676_), .B1(new_n790_), .B2(new_n802_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n810_), .ZN(G1341gat));
  NAND2_X1  g613(.A1(new_n790_), .A2(new_n802_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n323_), .A2(G127gat), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT121), .Z(new_n817_));
  OAI21_X1  g616(.A(new_n323_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n818_));
  INV_X1    g617(.A(G127gat), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n815_), .A2(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(G1342gat));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n785_), .A2(KEYINPUT119), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n800_), .A2(new_n804_), .A3(new_n729_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n688_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n821_), .B1(new_n824_), .B2(G134gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n598_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n826_));
  INV_X1    g625(.A(G134gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT122), .A3(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(G134gat), .B(new_n628_), .C1(new_n789_), .C2(new_n801_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n825_), .A2(new_n828_), .A3(new_n829_), .ZN(G1343gat));
  NAND2_X1  g629(.A1(new_n798_), .A2(new_n799_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(new_n595_), .A3(new_n526_), .A4(new_n613_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT123), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n806_), .A2(new_n474_), .A3(new_n540_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n526_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G141gat), .B1(new_n837_), .B2(new_n590_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n833_), .A2(new_n836_), .ZN(new_n839_));
  INV_X1    g638(.A(G141gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n589_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(G1344gat));
  OAI21_X1  g641(.A(G148gat), .B1(new_n837_), .B2(new_n676_), .ZN(new_n843_));
  INV_X1    g642(.A(G148gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n839_), .A2(new_n844_), .A3(new_n567_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1345gat));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n839_), .A2(new_n323_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n839_), .B2(new_n323_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1346gat));
  AOI21_X1  g649(.A(G162gat), .B1(new_n839_), .B2(new_n598_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n837_), .A2(new_n290_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(G162gat), .ZN(G1347gat));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n613_), .A2(new_n595_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n424_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n589_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT124), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n858_), .A2(KEYINPUT124), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n800_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT125), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(G169gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n861_), .B2(G169gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n854_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n865_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT62), .A3(new_n863_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n800_), .A2(new_n589_), .A3(new_n330_), .A4(new_n857_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n868_), .A3(new_n869_), .ZN(G1348gat));
  NAND2_X1  g669(.A1(new_n800_), .A2(new_n857_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n676_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n331_), .ZN(G1349gat));
  NOR2_X1   g672(.A1(new_n871_), .A2(new_n622_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(KEYINPUT126), .A3(G183gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n383_), .B1(new_n876_), .B2(new_n349_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n874_), .B2(new_n877_), .ZN(G1350gat));
  OAI21_X1  g677(.A(G190gat), .B1(new_n871_), .B2(new_n290_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n598_), .B1(new_n346_), .B2(new_n384_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n871_), .B2(new_n880_), .ZN(G1351gat));
  NOR3_X1   g680(.A1(new_n540_), .A2(new_n595_), .A3(new_n494_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n806_), .B1(KEYINPUT127), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT127), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n604_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n589_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n567_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g691(.A(KEYINPUT63), .B(G211gat), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n887_), .A2(new_n622_), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n888_), .A2(new_n323_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(G1354gat));
  NOR3_X1   g696(.A1(new_n887_), .A2(new_n364_), .A3(new_n290_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n888_), .A2(new_n598_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n364_), .B2(new_n899_), .ZN(G1355gat));
endmodule


