//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n967_, new_n968_, new_n969_, new_n970_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n984_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n992_, new_n993_;
  XOR2_X1   g000(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT25), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G190gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  OR3_X1    g022(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n218_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n213_), .A2(KEYINPUT81), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G176gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n212_), .A2(KEYINPUT22), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT82), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT81), .B(G176gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G169gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n233_), .A2(KEYINPUT83), .A3(new_n237_), .A4(new_n215_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT84), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n220_), .A2(new_n222_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n203_), .A2(new_n207_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n221_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n232_), .A2(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT83), .B1(new_n245_), .B2(new_n237_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n225_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G218gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G211gat), .ZN(new_n249_));
  INV_X1    g048(.A(G211gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G218gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n253_));
  INV_X1    g052(.A(G197gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT21), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(G197gat), .B2(G204gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n252_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n253_), .A2(G197gat), .A3(new_n255_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n254_), .A3(G204gat), .ZN(new_n262_));
  INV_X1    g061(.A(G204gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT91), .B1(new_n263_), .B2(G197gat), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n260_), .A2(new_n257_), .A3(new_n262_), .A4(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n257_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT92), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT92), .B1(new_n267_), .B2(new_n268_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n266_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n247_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT95), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n240_), .A2(new_n242_), .A3(new_n224_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n217_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n240_), .A2(KEYINPUT95), .A3(new_n242_), .A4(new_n224_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT96), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n235_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n235_), .A2(new_n279_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n234_), .A3(new_n281_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n223_), .A2(new_n241_), .B1(G169gat), .B2(G176gat), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n277_), .A2(new_n278_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n253_), .A2(G197gat), .A3(new_n255_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n264_), .A2(new_n262_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n268_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n289_), .A2(new_n269_), .B1(new_n265_), .B2(new_n259_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n274_), .B1(new_n284_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT19), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n273_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n276_), .A2(new_n275_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n218_), .A3(new_n278_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n282_), .A2(new_n283_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n274_), .B1(new_n272_), .B2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n290_), .B(new_n225_), .C1(new_n246_), .C2(new_n244_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n294_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT18), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G64gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G92gat), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n295_), .A2(new_n302_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n247_), .A2(new_n272_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT20), .B1(new_n284_), .B2(new_n290_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n293_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n273_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n308_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n202_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n300_), .A2(new_n301_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(new_n293_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n294_), .B1(new_n273_), .B2(new_n291_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n306_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n308_), .A3(new_n312_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT27), .A3(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n314_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322_));
  INV_X1    g121(.A(G141gat), .ZN(new_n323_));
  INV_X1    g122(.A(G148gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .A4(KEYINPUT89), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT89), .ZN(new_n326_));
  OAI22_X1  g125(.A1(new_n326_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n325_), .A2(new_n327_), .A3(new_n330_), .A4(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n337_), .A2(new_n328_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n333_), .A2(new_n340_), .A3(new_n334_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G120gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G113gat), .ZN(new_n345_));
  INV_X1    g144(.A(G113gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G120gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT86), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT86), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n345_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n351_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n350_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n343_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n332_), .A2(new_n335_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n355_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n352_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT97), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n357_), .A2(new_n353_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT97), .A3(new_n359_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n358_), .A2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n367_), .A2(G225gat), .A3(G233gat), .A4(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G1gat), .B(G29gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT0), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G57gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G85gat), .ZN(new_n375_));
  INV_X1    g174(.A(G57gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n373_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G85gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n364_), .A2(new_n382_), .A3(new_n366_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n370_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT98), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n370_), .A2(KEYINPUT98), .A3(new_n381_), .A4(new_n383_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n370_), .A2(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n380_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G22gat), .B(G50gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT28), .ZN(new_n393_));
  OR3_X1    g192(.A1(new_n343_), .A2(KEYINPUT29), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT94), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n343_), .B2(KEYINPUT29), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n395_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n289_), .A2(new_n269_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT93), .B1(new_n402_), .B2(new_n266_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n401_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n404_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n400_), .B(new_n406_), .C1(new_n290_), .C2(KEYINPUT93), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n272_), .B1(new_n408_), .B2(new_n359_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n399_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n405_), .A2(new_n407_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n409_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n398_), .A3(new_n410_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n321_), .A2(new_n391_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n247_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT30), .B(new_n225_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G15gat), .B(G43gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n365_), .B(KEYINPUT31), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n421_), .A2(new_n422_), .A3(new_n428_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n421_), .A2(new_n422_), .A3(new_n428_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n428_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(KEYINPUT85), .A3(new_n433_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n432_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n434_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI211_X1 g241(.A(KEYINPUT87), .B(new_n432_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n419_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n438_), .A2(new_n439_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT87), .B1(new_n448_), .B2(new_n432_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(new_n441_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(KEYINPUT88), .A4(new_n434_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n447_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n381_), .B1(new_n370_), .B2(new_n383_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n385_), .B2(new_n384_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT32), .ZN(new_n455_));
  OAI22_X1  g254(.A1(new_n295_), .A2(new_n302_), .B1(new_n455_), .B2(new_n306_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n317_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n306_), .A2(new_n455_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n457_), .B(new_n458_), .C1(new_n293_), .C2(new_n315_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n454_), .A2(new_n387_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n367_), .A2(new_n369_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n382_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n382_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n380_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n453_), .B2(KEYINPUT33), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n306_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n319_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469_));
  AOI211_X1 g268(.A(new_n469_), .B(new_n381_), .C1(new_n370_), .C2(new_n383_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n466_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n418_), .B1(new_n460_), .B2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n390_), .A2(new_n418_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT100), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n321_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n454_), .A2(new_n387_), .A3(new_n417_), .A4(new_n413_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n314_), .A2(new_n320_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT100), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n445_), .B1(new_n452_), .B2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G85gat), .B(G92gat), .Z(new_n481_));
  NOR2_X1   g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(KEYINPUT66), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  OAI22_X1  g284(.A1(new_n485_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n481_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT8), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT10), .B(G99gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT64), .B(G106gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n492_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G92gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT65), .B1(new_n378_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT9), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n378_), .A2(new_n499_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT9), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT65), .B(new_n503_), .C1(new_n378_), .C2(new_n499_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT8), .B(new_n481_), .C1(new_n487_), .C2(new_n492_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n495_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT12), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n376_), .A2(G64gat), .ZN(new_n512_));
  INV_X1    g311(.A(G64gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(G57gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(G57gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n376_), .A2(G64gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT67), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G71gat), .B(G78gat), .Z(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n515_), .A2(new_n519_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(KEYINPUT11), .ZN(new_n525_));
  AOI211_X1 g324(.A(KEYINPUT68), .B(new_n516_), .C1(new_n515_), .C2(new_n519_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT67), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT67), .B1(new_n517_), .B2(new_n518_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT11), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT68), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n523_), .A3(KEYINPUT11), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n527_), .A2(new_n533_), .A3(KEYINPUT70), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT70), .B1(new_n527_), .B2(new_n533_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n510_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n525_), .A2(new_n526_), .A3(new_n522_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n531_), .A2(new_n532_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n508_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n495_), .A2(new_n507_), .A3(new_n506_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n527_), .A3(new_n533_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT12), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n536_), .A2(KEYINPUT71), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n527_), .A2(new_n533_), .A3(KEYINPUT70), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n509_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n543_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n544_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT69), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G120gat), .B(G148gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n263_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT5), .B(G176gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n551_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(KEYINPUT13), .A3(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G169gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n254_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT76), .ZN(new_n570_));
  INV_X1    g369(.A(G1gat), .ZN(new_n571_));
  INV_X1    g370(.A(G8gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT75), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT75), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(G8gat), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT14), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n570_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT75), .B(G8gat), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT76), .B(KEYINPUT14), .C1(new_n579_), .C2(new_n571_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G15gat), .B(G22gat), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(G1gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n571_), .A3(new_n583_), .ZN(new_n586_));
  AOI21_X1  g385(.A(G8gat), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n571_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n588_));
  AOI211_X1 g387(.A(G1gat), .B(new_n582_), .C1(new_n578_), .C2(new_n580_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n572_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G29gat), .B(G36gat), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT72), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G36gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(G29gat), .ZN(new_n596_));
  INV_X1    g395(.A(G29gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G36gat), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n596_), .A2(new_n598_), .A3(new_n593_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G43gat), .B1(new_n594_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT72), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n592_), .A2(new_n593_), .ZN(new_n603_));
  INV_X1    g402(.A(G43gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(G50gat), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(G50gat), .A3(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n591_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n585_), .A2(G8gat), .A3(new_n586_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n572_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n610_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT79), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT79), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n617_), .B(new_n610_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n611_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT15), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n610_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n608_), .A2(KEYINPUT15), .A3(new_n609_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n591_), .A2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n620_), .B(KEYINPUT80), .Z(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n627_), .B(new_n629_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n569_), .B1(new_n622_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n614_), .A2(new_n615_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n615_), .B1(new_n587_), .B2(new_n590_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n617_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n614_), .A2(KEYINPUT79), .A3(new_n615_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n633_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n630_), .B(new_n569_), .C1(new_n637_), .C2(new_n620_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n480_), .A2(new_n566_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n591_), .B(new_n642_), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n643_), .A2(new_n538_), .A3(new_n537_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n538_), .B2(new_n537_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT78), .ZN(new_n647_));
  XOR2_X1   g446(.A(G127gat), .B(G155gat), .Z(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(G183gat), .B(G211gat), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT17), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n644_), .A2(new_n645_), .A3(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n534_), .A2(new_n535_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n643_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n643_), .A2(new_n654_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n655_), .A2(KEYINPUT17), .A3(new_n656_), .A4(new_n651_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G190gat), .B(G218gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(G134gat), .B(G162gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT36), .Z(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT74), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n626_), .A2(new_n508_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(G232gat), .A2(G233gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT34), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT35), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n615_), .A2(new_n540_), .B1(new_n668_), .B2(new_n667_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n664_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n664_), .B2(new_n671_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n663_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n674_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n661_), .A2(KEYINPUT36), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n672_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n663_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n676_), .B2(new_n672_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n679_), .B(KEYINPUT37), .C1(KEYINPUT73), .C2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT37), .B1(new_n681_), .B2(KEYINPUT73), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n675_), .A2(new_n678_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n658_), .B1(new_n682_), .B2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n641_), .A2(new_n571_), .A3(new_n390_), .A4(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n689_));
  OR2_X1    g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n658_), .A2(new_n684_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n641_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G1gat), .B1(new_n692_), .B2(new_n391_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n688_), .A2(new_n689_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n690_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT102), .ZN(G1324gat));
  OAI21_X1  g495(.A(G8gat), .B1(new_n692_), .B2(new_n321_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT39), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT39), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n641_), .A2(new_n686_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n477_), .A2(new_n579_), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n698_), .A2(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g502(.A(new_n452_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n641_), .A2(new_n704_), .A3(new_n691_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G15gat), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT103), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT103), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n709_));
  OR3_X1    g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n700_), .A2(G15gat), .A3(new_n452_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(G1326gat));
  OAI21_X1  g512(.A(G22gat), .B1(new_n692_), .B2(new_n418_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT42), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n418_), .A2(G22gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n700_), .B2(new_n716_), .ZN(G1327gat));
  INV_X1    g516(.A(new_n658_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(new_n679_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n641_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n597_), .A3(new_n390_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n682_), .A2(new_n685_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n480_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n480_), .C2(new_n723_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n480_), .A2(KEYINPUT43), .A3(new_n723_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n566_), .A2(new_n718_), .A3(new_n640_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT105), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n729_), .A2(new_n734_), .A3(new_n730_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n729_), .A2(KEYINPUT44), .A3(new_n730_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n390_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n597_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT106), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(KEYINPUT106), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n722_), .B1(new_n740_), .B2(new_n741_), .ZN(G1328gat));
  AND3_X1   g541(.A1(new_n729_), .A2(new_n734_), .A3(new_n730_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n734_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(KEYINPUT44), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n737_), .A2(new_n477_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G36gat), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n477_), .A2(new_n595_), .ZN(new_n751_));
  OR3_X1    g550(.A1(new_n720_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n720_), .B2(new_n751_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .A4(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n748_), .A2(new_n749_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n758_));
  INV_X1    g557(.A(new_n746_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n595_), .B1(new_n736_), .B2(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n757_), .B(new_n758_), .C1(new_n760_), .C2(new_n754_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n756_), .A2(new_n761_), .ZN(G1329gat));
  INV_X1    g561(.A(new_n444_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n737_), .A2(G43gat), .A3(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n745_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n721_), .A2(new_n704_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n604_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT108), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n765_), .A2(KEYINPUT47), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT47), .B1(new_n765_), .B2(new_n768_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1330gat));
  INV_X1    g570(.A(new_n418_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n737_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n607_), .B1(new_n736_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n418_), .A2(G50gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT109), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n720_), .A2(new_n777_), .ZN(new_n778_));
  OR3_X1    g577(.A1(new_n774_), .A2(new_n775_), .A3(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1331gat));
  NOR2_X1   g580(.A1(new_n480_), .A2(new_n639_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT112), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n686_), .A2(new_n566_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT111), .Z(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT113), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n390_), .A2(new_n376_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n782_), .A2(new_n566_), .A3(new_n691_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(new_n391_), .ZN(new_n791_));
  OAI22_X1  g590(.A1(new_n787_), .A2(new_n788_), .B1(new_n376_), .B2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT114), .ZN(G1332gat));
  AOI21_X1  g592(.A(new_n513_), .B1(new_n789_), .B2(new_n477_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT48), .Z(new_n795_));
  NAND2_X1  g594(.A1(new_n477_), .A2(new_n513_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n787_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT115), .ZN(G1333gat));
  INV_X1    g597(.A(G71gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n789_), .B2(new_n704_), .ZN(new_n800_));
  XOR2_X1   g599(.A(new_n800_), .B(KEYINPUT49), .Z(new_n801_));
  NAND2_X1  g600(.A1(new_n704_), .A2(new_n799_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n787_), .B2(new_n802_), .ZN(G1334gat));
  INV_X1    g602(.A(G78gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n789_), .B2(new_n772_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT50), .Z(new_n806_));
  NAND2_X1  g605(.A1(new_n772_), .A2(new_n804_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n787_), .B2(new_n807_), .ZN(G1335gat));
  NAND2_X1  g607(.A1(new_n566_), .A2(new_n658_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n639_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n729_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G85gat), .B1(new_n811_), .B2(new_n391_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n809_), .A2(new_n679_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n783_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n390_), .A2(new_n378_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n812_), .B1(new_n814_), .B2(new_n815_), .ZN(G1336gat));
  OAI21_X1  g615(.A(G92gat), .B1(new_n811_), .B2(new_n321_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n477_), .A2(new_n499_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n814_), .B2(new_n818_), .ZN(G1337gat));
  OR2_X1    g618(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n729_), .A2(new_n704_), .A3(new_n810_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n821_), .A2(KEYINPUT116), .A3(G99gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT116), .B1(new_n821_), .B2(G99gat), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n814_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n763_), .A2(new_n496_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n825_), .A2(new_n826_), .B1(KEYINPUT117), .B2(KEYINPUT51), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n820_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n827_), .B(new_n820_), .C1(new_n823_), .C2(new_n822_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1338gat));
  NAND3_X1  g630(.A1(new_n825_), .A2(new_n497_), .A3(new_n772_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n729_), .A2(new_n772_), .A3(new_n810_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n833_), .A2(new_n834_), .A3(G106gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n833_), .B2(G106gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT58), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n627_), .B(new_n628_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n569_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(new_n842_), .C1(new_n637_), .C2(new_n628_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n561_), .A2(new_n638_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n544_), .B1(new_n543_), .B2(new_n550_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n551_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n542_), .A2(new_n539_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n849_));
  AOI211_X1 g648(.A(KEYINPUT71), .B(new_n509_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n544_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n846_), .A4(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n558_), .B1(new_n847_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n844_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT56), .B(new_n558_), .C1(new_n847_), .C2(new_n853_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n840_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n849_), .A2(new_n851_), .A3(new_n850_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n851_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(KEYINPUT55), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n559_), .B1(new_n861_), .B2(new_n852_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT56), .ZN(new_n863_));
  INV_X1    g662(.A(new_n840_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n854_), .A2(new_n855_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .A4(new_n844_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n723_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n858_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n862_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n854_), .A2(new_n869_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n638_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n561_), .B1(new_n873_), .B2(new_n631_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(new_n872_), .A3(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n562_), .A2(new_n638_), .A3(new_n843_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n684_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n868_), .B1(new_n878_), .B2(KEYINPUT57), .ZN(new_n879_));
  INV_X1    g678(.A(new_n877_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n874_), .B1(new_n854_), .B2(new_n869_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n871_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n882_), .A2(new_n883_), .A3(new_n684_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n658_), .B1(new_n879_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n566_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n639_), .B1(KEYINPUT118), .B2(KEYINPUT54), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n686_), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n890_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n886_), .A2(new_n686_), .A3(new_n887_), .A4(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n885_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n418_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n477_), .A2(new_n391_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n444_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(new_n346_), .A3(new_n639_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n772_), .B1(new_n885_), .B2(new_n895_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n900_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n883_), .B1(new_n882_), .B2(new_n684_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n876_), .A2(new_n877_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(KEYINPUT57), .A3(new_n679_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n909_), .A3(new_n868_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n894_), .B1(new_n910_), .B2(new_n658_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n911_), .A2(KEYINPUT59), .A3(new_n772_), .A4(new_n901_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n906_), .A2(new_n912_), .A3(new_n640_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n903_), .B1(new_n913_), .B2(new_n346_), .ZN(G1340gat));
  NOR2_X1   g713(.A1(new_n886_), .A2(G120gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n902_), .B1(KEYINPUT60), .B2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n906_), .A2(new_n912_), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n916_), .A2(new_n566_), .A3(new_n917_), .ZN(new_n918_));
  OAI22_X1  g717(.A1(new_n918_), .A2(new_n344_), .B1(KEYINPUT60), .B2(new_n916_), .ZN(G1341gat));
  AOI21_X1  g718(.A(G127gat), .B1(new_n902_), .B2(new_n718_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT121), .B(G127gat), .Z(new_n921_));
  NAND2_X1  g720(.A1(new_n718_), .A2(new_n921_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(KEYINPUT122), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n920_), .B1(new_n917_), .B2(new_n923_), .ZN(G1342gat));
  INV_X1    g723(.A(G134gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n917_), .B2(new_n867_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n902_), .A2(new_n925_), .A3(new_n684_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT123), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n906_), .A2(new_n912_), .A3(new_n723_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n930_), .B(new_n927_), .C1(new_n931_), .C2(new_n925_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n932_), .ZN(G1343gat));
  NAND4_X1  g732(.A1(new_n896_), .A2(new_n452_), .A3(new_n772_), .A4(new_n898_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n639_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G141gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n936_), .A2(new_n323_), .A3(new_n639_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1344gat));
  XOR2_X1   g739(.A(KEYINPUT125), .B(G148gat), .Z(new_n941_));
  AND3_X1   g740(.A1(new_n936_), .A2(new_n566_), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n936_), .B2(new_n566_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1345gat));
  NAND2_X1  g743(.A1(new_n936_), .A2(new_n718_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT61), .B(G155gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n946_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n936_), .A2(new_n718_), .A3(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1346gat));
  NAND2_X1  g749(.A1(new_n936_), .A2(new_n684_), .ZN(new_n951_));
  INV_X1    g750(.A(G162gat), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n867_), .A2(G162gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT126), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n951_), .A2(new_n952_), .B1(new_n936_), .B2(new_n954_), .ZN(G1347gat));
  NAND3_X1  g754(.A1(new_n704_), .A2(new_n391_), .A3(new_n477_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n897_), .A2(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n212_), .B1(new_n957_), .B2(new_n639_), .ZN(new_n958_));
  OR2_X1    g757(.A1(new_n958_), .A2(KEYINPUT62), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(KEYINPUT62), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n280_), .A2(new_n281_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n957_), .A2(new_n639_), .ZN(new_n962_));
  OAI211_X1 g761(.A(new_n959_), .B(new_n960_), .C1(new_n961_), .C2(new_n962_), .ZN(G1348gat));
  NAND2_X1  g762(.A1(new_n957_), .A2(new_n566_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n213_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n234_), .B2(new_n964_), .ZN(G1349gat));
  INV_X1    g765(.A(new_n957_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n967_), .A2(new_n658_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n968_), .A2(G183gat), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n204_), .A2(new_n206_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n969_), .B1(new_n968_), .B2(new_n970_), .ZN(G1350gat));
  OAI21_X1  g770(.A(G190gat), .B1(new_n967_), .B2(new_n723_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n684_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n967_), .B2(new_n973_), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n911_), .A2(new_n704_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n321_), .A2(new_n476_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  INV_X1    g776(.A(new_n977_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n978_), .A2(G197gat), .A3(new_n639_), .ZN(new_n979_));
  AND2_X1   g778(.A1(new_n979_), .A2(KEYINPUT127), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n979_), .A2(KEYINPUT127), .ZN(new_n981_));
  AOI21_X1  g780(.A(G197gat), .B1(new_n978_), .B2(new_n639_), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n980_), .A2(new_n981_), .A3(new_n982_), .ZN(G1352gat));
  NAND2_X1  g782(.A1(new_n978_), .A2(new_n566_), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n984_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n985_));
  AOI21_X1  g784(.A(new_n985_), .B1(new_n263_), .B2(new_n984_), .ZN(G1353gat));
  NAND2_X1  g785(.A1(new_n978_), .A2(new_n718_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n988_));
  AND2_X1   g787(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n989_));
  NOR3_X1   g788(.A1(new_n987_), .A2(new_n988_), .A3(new_n989_), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n990_), .B1(new_n987_), .B2(new_n988_), .ZN(G1354gat));
  OAI21_X1  g790(.A(G218gat), .B1(new_n977_), .B2(new_n723_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n684_), .A2(new_n248_), .ZN(new_n993_));
  OAI21_X1  g792(.A(new_n992_), .B1(new_n977_), .B2(new_n993_), .ZN(G1355gat));
endmodule


