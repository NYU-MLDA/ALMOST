//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_;
  INV_X1    g000(.A(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT66), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT7), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT67), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n207_), .B(new_n209_), .C1(new_n210_), .C2(new_n205_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT64), .B(G85gat), .Z(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n212_), .A4(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n221_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n203_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n223_), .A2(new_n224_), .A3(new_n209_), .A4(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n214_), .A2(new_n215_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n216_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G57gat), .B(G64gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G71gat), .B(G78gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n230_), .B(KEYINPUT11), .Z(new_n234_));
  OAI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(new_n232_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(KEYINPUT12), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT12), .B1(new_n236_), .B2(new_n237_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n235_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n216_), .A2(new_n240_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G230gat), .A2(G233gat), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n241_), .A2(KEYINPUT69), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT69), .B1(new_n241_), .B2(new_n242_), .ZN(new_n244_));
  OAI22_X1  g043(.A1(new_n238_), .A2(new_n239_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n236_), .A2(new_n241_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(G230gat), .A3(G233gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT5), .B(G176gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G204gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G120gat), .B(G148gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n250_), .B(new_n251_), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n252_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n245_), .A2(new_n247_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT13), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(KEYINPUT13), .A3(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G15gat), .B(G22gat), .ZN(new_n261_));
  INV_X1    g060(.A(G1gat), .ZN(new_n262_));
  INV_X1    g061(.A(G8gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT14), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G1gat), .B(G8gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G29gat), .B(G36gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G43gat), .B(G50gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n267_), .B(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n267_), .A2(new_n270_), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n270_), .B(KEYINPUT15), .Z(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(new_n267_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G229gat), .A2(G233gat), .ZN(new_n275_));
  MUX2_X1   g074(.A(new_n271_), .B(new_n274_), .S(new_n275_), .Z(new_n276_));
  XNOR2_X1  g075(.A(G113gat), .B(G141gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT78), .ZN(new_n278_));
  XOR2_X1   g077(.A(G169gat), .B(G197gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n276_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n260_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT98), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT97), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT23), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(G183gat), .A3(G190gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT24), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(KEYINPUT80), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n299_));
  INV_X1    g098(.A(new_n293_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n301_), .B2(new_n296_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT26), .B(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n295_), .A2(KEYINPUT24), .A3(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n298_), .A2(new_n302_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G176gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n310_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT22), .B(G169gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(KEYINPUT81), .A3(new_n310_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n316_), .A2(new_n318_), .A3(new_n306_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n287_), .A2(new_n293_), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  INV_X1    g120(.A(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT82), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n320_), .A2(KEYINPUT82), .A3(new_n323_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n319_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n309_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n328_));
  AND2_X1   g127(.A1(G211gat), .A2(G218gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G211gat), .A2(G218gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G197gat), .B(G204gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(KEYINPUT90), .ZN(new_n333_));
  INV_X1    g132(.A(G204gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G197gat), .ZN(new_n335_));
  INV_X1    g134(.A(G197gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G204gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n337_), .A3(KEYINPUT90), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT21), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n328_), .B1(new_n333_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT21), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n332_), .B2(KEYINPUT90), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n337_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT90), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n342_), .A2(KEYINPUT91), .A3(new_n345_), .A4(new_n331_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n335_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n341_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n331_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT92), .B1(new_n347_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT92), .ZN(new_n353_));
  AOI211_X1 g152(.A(new_n353_), .B(new_n350_), .C1(new_n340_), .C2(new_n346_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n327_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT20), .ZN(new_n356_));
  AND4_X1   g155(.A1(new_n320_), .A2(new_n305_), .A3(new_n297_), .A4(new_n307_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n317_), .A2(KEYINPUT94), .ZN(new_n358_));
  INV_X1    g157(.A(new_n313_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT94), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n311_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n294_), .A2(new_n323_), .B1(new_n362_), .B2(new_n310_), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n306_), .B(KEYINPUT93), .Z(new_n364_));
  AOI21_X1  g163(.A(new_n357_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n350_), .B1(new_n340_), .B2(new_n346_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n356_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n355_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT19), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n285_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  AOI211_X1 g171(.A(KEYINPUT97), .B(new_n372_), .C1(new_n355_), .C2(new_n367_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n347_), .A2(new_n351_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n353_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n366_), .A2(KEYINPUT92), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n326_), .A4(new_n309_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n294_), .A2(new_n323_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(new_n310_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(new_n364_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n357_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n356_), .B1(new_n382_), .B2(new_n374_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n377_), .A2(new_n372_), .A3(new_n383_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n371_), .A2(new_n373_), .A3(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(new_n219_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT18), .B(G64gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n284_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n368_), .A2(new_n370_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n372_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n391_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G113gat), .B(G120gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  INV_X1    g198(.A(G155gat), .ZN(new_n400_));
  INV_X1    g199(.A(G162gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT1), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT1), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G155gat), .A3(G162gat), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n402_), .B(new_n404_), .C1(G155gat), .C2(G162gat), .ZN(new_n405_));
  INV_X1    g204(.A(G141gat), .ZN(new_n406_));
  INV_X1    g205(.A(G148gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n405_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n400_), .A2(new_n401_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G155gat), .A2(G162gat), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT2), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n409_), .B1(new_n414_), .B2(KEYINPUT87), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n416_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n406_), .A2(new_n407_), .A3(KEYINPUT3), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(G141gat), .B2(G148gat), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n420_), .A2(new_n422_), .B1(KEYINPUT87), .B2(new_n414_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n413_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n399_), .B1(new_n410_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n413_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n420_), .A2(new_n422_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n414_), .A2(KEYINPUT87), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n429_), .B2(new_n418_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n397_), .B(new_n398_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n405_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n425_), .A2(new_n433_), .A3(KEYINPUT4), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n425_), .A2(KEYINPUT4), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n425_), .A2(new_n433_), .A3(KEYINPUT95), .A4(KEYINPUT4), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n425_), .A2(new_n433_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n437_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G57gat), .B(G85gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n447_), .B(new_n448_), .Z(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n441_), .A2(new_n443_), .A3(new_n449_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n396_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n355_), .A2(new_n367_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT97), .B1(new_n454_), .B2(new_n372_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n384_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n368_), .A2(new_n285_), .A3(new_n370_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(KEYINPUT98), .A3(new_n395_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n392_), .A2(new_n453_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT99), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n430_), .A2(new_n462_), .A3(new_n432_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G78gat), .B(G106gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G22gat), .B(G50gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n462_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G228gat), .A2(G233gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n472_), .B(KEYINPUT89), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n469_), .A2(new_n366_), .A3(new_n473_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n480_), .A3(new_n476_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n468_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n483_));
  AOI211_X1 g282(.A(new_n478_), .B(new_n475_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n467_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n466_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n481_), .A3(new_n468_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n467_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n465_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n452_), .A2(KEYINPUT33), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n441_), .A2(new_n443_), .A3(new_n491_), .A4(new_n449_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n454_), .A2(new_n372_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n377_), .A2(new_n383_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n494_), .B(new_n390_), .C1(new_n372_), .C2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n389_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n436_), .A2(new_n437_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n442_), .A2(new_n438_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n450_), .A3(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n493_), .A2(new_n496_), .A3(new_n497_), .A4(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n486_), .A2(new_n489_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT99), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n392_), .A2(new_n453_), .A3(new_n459_), .A4(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n461_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT30), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n327_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n327_), .B(KEYINPUT30), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G227gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT83), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G43gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n511_), .A2(new_n513_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n506_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n431_), .B(KEYINPUT31), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n511_), .A2(new_n513_), .A3(new_n519_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(KEYINPUT86), .A3(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n505_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n486_), .A2(new_n489_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n451_), .A2(new_n452_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT27), .ZN(new_n537_));
  INV_X1    g336(.A(new_n496_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n458_), .A2(new_n389_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n539_), .B2(KEYINPUT100), .ZN(new_n540_));
  OR3_X1    g339(.A1(new_n385_), .A2(KEYINPUT100), .A3(new_n390_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n537_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n496_), .A2(new_n537_), .A3(new_n497_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n536_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n530_), .A2(new_n533_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n531_), .A2(new_n534_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n283_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n229_), .A2(new_n270_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n229_), .A2(new_n273_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n549_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n550_), .A2(KEYINPUT72), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n553_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT71), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n555_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT36), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n558_), .B1(new_n550_), .B2(KEYINPUT72), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n565_), .A2(new_n550_), .A3(new_n554_), .A4(new_n549_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n559_), .A2(new_n566_), .B1(new_n569_), .B2(new_n562_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n548_), .B(KEYINPUT37), .C1(new_n568_), .C2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n559_), .A2(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n562_), .A2(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n567_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n267_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n240_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT75), .ZN(new_n582_));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT76), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n582_), .A2(new_n590_), .ZN(new_n591_));
  OR3_X1    g390(.A1(new_n581_), .A2(new_n588_), .A3(new_n587_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT77), .Z(new_n594_));
  NOR2_X1   g393(.A1(new_n578_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n547_), .A2(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n596_), .A2(G1gat), .A3(new_n536_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT38), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT101), .ZN(new_n599_));
  INV_X1    g398(.A(new_n546_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n574_), .A2(new_n567_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n593_), .A3(new_n283_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G1gat), .B1(new_n603_), .B2(new_n536_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n599_), .B(new_n604_), .C1(KEYINPUT38), .C2(new_n597_), .ZN(G1324gat));
  NOR2_X1   g404(.A1(new_n542_), .A2(new_n543_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G8gat), .B1(new_n603_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT39), .ZN(new_n609_));
  INV_X1    g408(.A(new_n596_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n263_), .A3(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(G1325gat));
  OAI21_X1  g413(.A(G15gat), .B1(new_n603_), .B2(new_n530_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT103), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT41), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n610_), .A2(new_n532_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(G15gat), .B2(new_n618_), .ZN(G1326gat));
  OAI21_X1  g418(.A(G22gat), .B1(new_n603_), .B2(new_n533_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n533_), .A2(G22gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n596_), .B2(new_n622_), .ZN(G1327gat));
  NAND2_X1  g422(.A1(new_n594_), .A2(new_n601_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT107), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n547_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G29gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n535_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n531_), .A2(new_n534_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n544_), .A2(new_n545_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n578_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n578_), .A3(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT43), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n546_), .A2(KEYINPUT104), .A3(new_n631_), .A4(new_n578_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n594_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n260_), .A2(new_n640_), .A3(new_n282_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n639_), .A2(new_n641_), .A3(KEYINPUT105), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT106), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n646_), .A2(new_n650_), .A3(new_n643_), .A4(new_n647_), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n536_), .B(new_n644_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n629_), .B1(new_n652_), .B2(new_n628_), .ZN(G1328gat));
  NOR3_X1   g452(.A1(new_n626_), .A2(G36gat), .A3(new_n607_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT45), .Z(new_n655_));
  INV_X1    g454(.A(KEYINPUT108), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n649_), .A2(new_n651_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n644_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n606_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n657_), .B1(new_n660_), .B2(G36gat), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(KEYINPUT108), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n661_), .B(new_n663_), .ZN(G1329gat));
  XNOR2_X1  g463(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n665_));
  OAI211_X1 g464(.A(G43gat), .B(new_n532_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT109), .B1(new_n658_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n669_));
  AOI211_X1 g468(.A(new_n669_), .B(new_n666_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G43gat), .B1(new_n627_), .B2(new_n532_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n665_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n665_), .ZN(new_n675_));
  NOR4_X1   g474(.A1(new_n668_), .A2(new_n670_), .A3(new_n672_), .A4(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1330gat));
  INV_X1    g476(.A(G50gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n533_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n627_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  AOI211_X1 g479(.A(new_n533_), .B(new_n644_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n678_), .ZN(G1331gat));
  NAND2_X1  g481(.A1(new_n595_), .A2(new_n260_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT111), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n600_), .A2(new_n281_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(KEYINPUT111), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n535_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n260_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n281_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n602_), .A2(new_n640_), .A3(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(new_n535_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n689_), .B1(G57gat), .B2(new_n693_), .ZN(G1332gat));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n606_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G64gat), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT48), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n607_), .A2(G64gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n687_), .B2(new_n698_), .ZN(G1333gat));
  INV_X1    g498(.A(G71gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n692_), .B2(new_n532_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT49), .Z(new_n702_));
  NAND3_X1  g501(.A1(new_n688_), .A2(new_n700_), .A3(new_n532_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1334gat));
  NAND2_X1  g503(.A1(new_n692_), .A2(new_n679_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G78gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT50), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n533_), .A2(G78gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n687_), .B2(new_n708_), .ZN(G1335gat));
  NAND3_X1  g508(.A1(new_n625_), .A2(new_n546_), .A3(new_n691_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT112), .ZN(new_n711_));
  AOI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n535_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n639_), .A2(new_n594_), .A3(new_n691_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n536_), .A2(new_n218_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(G1336gat));
  AOI21_X1  g514(.A(G92gat), .B1(new_n711_), .B2(new_n606_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n606_), .A2(G92gat), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT113), .Z(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n713_), .B2(new_n718_), .ZN(G1337gat));
  NAND3_X1  g518(.A1(new_n711_), .A2(new_n225_), .A3(new_n532_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT114), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT51), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n713_), .A2(new_n532_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n720_), .B(new_n722_), .C1(new_n202_), .C2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n721_), .A2(KEYINPUT51), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n724_), .B(new_n725_), .Z(G1338gat));
  NAND2_X1  g525(.A1(new_n713_), .A2(new_n679_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G106gat), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(KEYINPUT116), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(KEYINPUT116), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n731_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n711_), .A2(new_n203_), .A3(new_n679_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT53), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT53), .ZN(new_n738_));
  INV_X1    g537(.A(new_n733_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n730_), .A2(new_n731_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n738_), .B(new_n735_), .C1(new_n741_), .C2(new_n729_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n742_), .ZN(G1339gat));
  NAND3_X1  g542(.A1(new_n595_), .A2(new_n690_), .A3(new_n282_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT54), .Z(new_n745_));
  INV_X1    g544(.A(new_n593_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n255_), .A2(new_n281_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n241_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(G230gat), .A3(G233gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n245_), .A2(new_n752_), .ZN(new_n753_));
  OAI221_X1 g552(.A(KEYINPUT55), .B1(new_n243_), .B2(new_n244_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(KEYINPUT56), .A3(new_n252_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT56), .B1(new_n755_), .B2(new_n252_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n749_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n271_), .A2(new_n275_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n274_), .B(KEYINPUT118), .Z(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n275_), .ZN(new_n762_));
  MUX2_X1   g561(.A(new_n276_), .B(new_n762_), .S(new_n280_), .Z(new_n763_));
  AND3_X1   g562(.A1(new_n256_), .A2(KEYINPUT119), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT119), .B1(new_n256_), .B2(new_n763_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n759_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n601_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(KEYINPUT57), .A3(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n755_), .A2(new_n252_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n756_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n255_), .A3(new_n763_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n776_), .A2(KEYINPUT58), .A3(new_n255_), .A4(new_n763_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n578_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n771_), .A2(new_n772_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n745_), .B1(new_n746_), .B2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n606_), .A2(new_n536_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n533_), .A3(new_n532_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT120), .Z(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n281_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT121), .Z(new_n790_));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT57), .B1(new_n767_), .B2(new_n768_), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n770_), .B(new_n601_), .C1(new_n759_), .C2(new_n766_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n640_), .B1(new_n794_), .B2(new_n781_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n791_), .B(new_n786_), .C1(new_n795_), .C2(new_n745_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT122), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT59), .B1(new_n783_), .B2(new_n787_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n782_), .A2(new_n594_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n745_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT122), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n791_), .A4(new_n786_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n797_), .A2(new_n798_), .A3(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n281_), .A2(G113gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n790_), .B1(new_n804_), .B2(new_n805_), .ZN(G1340gat));
  NAND4_X1  g605(.A1(new_n797_), .A2(new_n260_), .A3(new_n798_), .A4(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G120gat), .ZN(new_n808_));
  INV_X1    g607(.A(G120gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n690_), .B2(KEYINPUT60), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n788_), .B(new_n810_), .C1(KEYINPUT60), .C2(new_n809_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT123), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n808_), .A2(KEYINPUT123), .A3(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1341gat));
  AOI21_X1  g615(.A(G127gat), .B1(new_n788_), .B2(new_n640_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n804_), .A2(G127gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n593_), .ZN(G1342gat));
  AOI21_X1  g618(.A(G134gat), .B1(new_n788_), .B2(new_n601_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n804_), .A2(new_n578_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g621(.A1(new_n607_), .A2(new_n535_), .ZN(new_n823_));
  NOR4_X1   g622(.A1(new_n783_), .A2(new_n533_), .A3(new_n532_), .A4(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n281_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n260_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n640_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G155gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n824_), .A2(new_n400_), .A3(new_n640_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n832_), .B(new_n834_), .ZN(G1346gat));
  AOI21_X1  g634(.A(G162gat), .B1(new_n824_), .B2(new_n601_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n578_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n401_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n824_), .B2(new_n838_), .ZN(G1347gat));
  NOR2_X1   g638(.A1(new_n607_), .A2(new_n535_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n534_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n801_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(G169gat), .B1(new_n843_), .B2(new_n282_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT62), .ZN(new_n845_));
  INV_X1    g644(.A(new_n843_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n281_), .A3(new_n362_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1348gat));
  AOI21_X1  g647(.A(G176gat), .B1(new_n846_), .B2(new_n260_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n783_), .A2(new_n534_), .A3(new_n841_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n690_), .A2(new_n310_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(G1349gat));
  AOI21_X1  g651(.A(G183gat), .B1(new_n850_), .B2(new_n640_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n843_), .A2(new_n746_), .A3(new_n303_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n843_), .B2(new_n837_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT125), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n846_), .A2(new_n601_), .A3(new_n304_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1351gat));
  NOR4_X1   g658(.A1(new_n783_), .A2(new_n533_), .A3(new_n532_), .A4(new_n841_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n281_), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n861_), .A2(KEYINPUT126), .A3(new_n336_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n336_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT126), .B1(new_n861_), .B2(new_n336_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(G1352gat));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n260_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n866_), .B(new_n867_), .Z(G1353gat));
  AND2_X1   g667(.A1(new_n860_), .A2(new_n593_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n869_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT63), .B(G211gat), .Z(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(new_n871_), .ZN(G1354gat));
  AOI21_X1  g671(.A(G218gat), .B1(new_n860_), .B2(new_n601_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n578_), .A2(G218gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n860_), .B2(new_n874_), .ZN(G1355gat));
endmodule


