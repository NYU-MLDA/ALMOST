//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(KEYINPUT84), .A3(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT84), .B1(new_n204_), .B2(G197gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT21), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n207_), .B(KEYINPUT85), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(new_n206_), .B2(G204gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n210_), .B(new_n211_), .C1(new_n213_), .C2(KEYINPUT21), .ZN(new_n214_));
  INV_X1    g013(.A(new_n211_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(KEYINPUT21), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT86), .B1(new_n214_), .B2(new_n216_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n227_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT77), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT23), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n224_), .A2(KEYINPUT24), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT78), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n236_), .B1(G183gat), .B2(G190gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT22), .B(G169gat), .Z(new_n242_));
  OAI211_X1 g041(.A(new_n241_), .B(new_n225_), .C1(G176gat), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n203_), .B1(new_n221_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G226gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT19), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n238_), .A2(new_n231_), .A3(new_n226_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n245_), .B(new_n248_), .C1(new_n217_), .C2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n217_), .A2(new_n250_), .ZN(new_n252_));
  OAI211_X1 g051(.A(KEYINPUT20), .B(new_n252_), .C1(new_n221_), .C2(new_n244_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n247_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G8gat), .B(G36gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(G64gat), .B(G92gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n255_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n217_), .B(KEYINPUT88), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n245_), .B1(new_n268_), .B2(new_n250_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n247_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n263_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(new_n262_), .A3(KEYINPUT27), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n267_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G78gat), .B(G106gat), .ZN(new_n275_));
  INV_X1    g074(.A(G228gat), .ZN(new_n276_));
  INV_X1    g075(.A(G233gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT83), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT3), .ZN(new_n284_));
  OR3_X1    g083(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n284_), .A2(new_n285_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n282_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(KEYINPUT1), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n283_), .B(new_n286_), .C1(new_n281_), .C2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT29), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n279_), .B1(new_n268_), .B2(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n279_), .B(new_n296_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n275_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n295_), .A2(KEYINPUT29), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G22gat), .B(G50gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT28), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n303_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n275_), .B(KEYINPUT89), .Z(new_n308_));
  NOR3_X1   g107(.A1(new_n299_), .A2(new_n301_), .A3(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT90), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n306_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n268_), .A2(new_n298_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n278_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n314_), .B2(new_n300_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n311_), .B1(new_n315_), .B2(new_n309_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n312_), .A3(new_n300_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n317_), .A2(new_n302_), .A3(new_n318_), .A4(new_n306_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n310_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT91), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n310_), .A2(KEYINPUT91), .A3(new_n316_), .A4(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n244_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G15gat), .B(G43gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT81), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT30), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n333_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(KEYINPUT82), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341_));
  INV_X1    g140(.A(G113gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G120gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT31), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n337_), .A2(KEYINPUT82), .A3(new_n339_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT82), .B1(new_n337_), .B2(new_n339_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n350_), .B2(new_n346_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n324_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n322_), .A2(new_n351_), .A3(new_n323_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n274_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n344_), .B(new_n295_), .Z(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT4), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(KEYINPUT93), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n344_), .A2(new_n295_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n358_), .B(new_n361_), .C1(KEYINPUT4), .C2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G1gat), .B(G29gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n356_), .B1(new_n365_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n363_), .A2(new_n364_), .A3(new_n370_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n373_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n324_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n271_), .A2(KEYINPUT32), .A3(new_n261_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT32), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n256_), .B1(new_n379_), .B2(new_n263_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n374_), .A2(new_n378_), .A3(new_n375_), .A4(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n373_), .B(KEYINPUT33), .ZN(new_n382_));
  INV_X1    g181(.A(new_n359_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n358_), .B1(KEYINPUT4), .B2(new_n362_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n357_), .B(KEYINPUT95), .Z(new_n385_));
  OAI221_X1 g184(.A(new_n371_), .B1(new_n383_), .B2(new_n384_), .C1(new_n385_), .C2(new_n360_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n382_), .A2(new_n262_), .A3(new_n264_), .A4(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n351_), .B1(new_n381_), .B2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n355_), .A2(new_n376_), .B1(new_n377_), .B2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G113gat), .B(G141gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(new_n222_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(new_n206_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G29gat), .B(G36gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G43gat), .ZN(new_n394_));
  INV_X1    g193(.A(G50gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n393_), .A2(G43gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(G43gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(G50gat), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G22gat), .ZN(new_n401_));
  INV_X1    g200(.A(G1gat), .ZN(new_n402_));
  INV_X1    g201(.A(G8gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT14), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G8gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT15), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT69), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n396_), .A2(new_n410_), .A3(new_n399_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(KEYINPUT15), .A3(new_n411_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n408_), .B1(new_n417_), .B2(new_n407_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G229gat), .A2(G233gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT75), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT75), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n400_), .B(new_n407_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n419_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n392_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n392_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n418_), .A2(new_n419_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n420_), .B(new_n428_), .C1(new_n429_), .C2(new_n425_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n202_), .B1(new_n389_), .B2(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n267_), .A2(new_n273_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n354_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n351_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n434_), .B(new_n376_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n388_), .A2(new_n377_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(KEYINPUT98), .A3(new_n431_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n433_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT7), .ZN(new_n442_));
  INV_X1    g241(.A(G99gat), .ZN(new_n443_));
  INV_X1    g242(.A(G106gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G99gat), .A2(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(G85gat), .A2(G92gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT65), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n443_), .A2(KEYINPUT10), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT10), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(G99gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(G106gat), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n448_), .A2(new_n449_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT9), .B1(new_n452_), .B2(new_n453_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(KEYINPUT64), .A3(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT64), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n464_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n451_), .A2(KEYINPUT65), .A3(new_n454_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT8), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT65), .B1(new_n451_), .B2(new_n454_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n458_), .B(new_n472_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(G57gat), .A2(G64gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G57gat), .A2(G64gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT11), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G57gat), .ZN(new_n480_));
  INV_X1    g279(.A(G64gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT11), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G57gat), .A2(G64gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(G78gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G71gat), .ZN(new_n487_));
  INV_X1    g286(.A(G71gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G78gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n479_), .A2(new_n485_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n482_), .A2(new_n484_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(KEYINPUT11), .A3(new_n487_), .A4(new_n489_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n491_), .A2(KEYINPUT66), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT66), .B1(new_n491_), .B2(new_n493_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n476_), .A2(new_n496_), .A3(KEYINPUT12), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n462_), .A2(new_n463_), .A3(new_n470_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n457_), .A2(new_n475_), .B1(new_n498_), .B2(new_n469_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n455_), .A2(new_n456_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(KEYINPUT8), .A3(new_n473_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n491_), .A2(new_n493_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n499_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G230gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n502_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT12), .B1(new_n476_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n504_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n476_), .A2(new_n506_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n503_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n505_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G120gat), .B(G148gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(new_n204_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT5), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(new_n223_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n509_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT13), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(KEYINPUT13), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT67), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(KEYINPUT67), .A3(new_n524_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT68), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(KEYINPUT73), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n407_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(new_n502_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT16), .B(G183gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G211gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n534_), .B1(KEYINPUT17), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(KEYINPUT17), .B2(new_n538_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n533_), .B(new_n496_), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(KEYINPUT17), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT74), .Z(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT37), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT15), .B1(new_n415_), .B2(new_n411_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n412_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n476_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT34), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT35), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI22_X1  g353(.A1(new_n476_), .A2(new_n400_), .B1(KEYINPUT35), .B2(new_n551_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n549_), .A2(KEYINPUT70), .A3(new_n554_), .A4(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(KEYINPUT70), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n554_), .A2(KEYINPUT70), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n474_), .A2(new_n475_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n458_), .A2(new_n472_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n558_), .B(new_n559_), .C1(new_n563_), .C2(new_n555_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT71), .B(G134gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n557_), .A2(new_n564_), .A3(KEYINPUT36), .A4(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT72), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n557_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n568_), .A2(KEYINPUT36), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n569_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n571_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n546_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n569_), .A2(new_n572_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n571_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(KEYINPUT37), .A3(new_n573_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n545_), .B1(new_n576_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n530_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n441_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n376_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(KEYINPUT38), .A3(new_n402_), .A4(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n441_), .A2(new_n585_), .A3(new_n583_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n590_), .A2(KEYINPUT99), .A3(KEYINPUT38), .A4(new_n402_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n529_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n431_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT100), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n574_), .A2(new_n575_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(new_n545_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n598_), .A3(new_n439_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT101), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n376_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n601_), .A2(KEYINPUT38), .B1(new_n402_), .B2(new_n590_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT102), .B1(new_n592_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(KEYINPUT38), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n590_), .A2(new_n402_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n606_), .A2(new_n607_), .A3(new_n588_), .A4(new_n591_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n608_), .ZN(G1324gat));
  OAI21_X1  g408(.A(G8gat), .B1(new_n599_), .B2(new_n434_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT39), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n434_), .A2(G8gat), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n584_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n612_), .B1(new_n584_), .B2(new_n613_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT40), .B(new_n611_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n600_), .B2(new_n352_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT41), .ZN(new_n622_));
  INV_X1    g421(.A(new_n584_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n623_), .A2(G15gat), .A3(new_n352_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n622_), .A2(new_n624_), .ZN(G1326gat));
  OAI21_X1  g424(.A(G22gat), .B1(new_n600_), .B2(new_n377_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT42), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n377_), .A2(G22gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n623_), .B2(new_n628_), .ZN(G1327gat));
  XNOR2_X1  g428(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n576_), .A2(new_n580_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n630_), .B1(new_n389_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633_));
  INV_X1    g432(.A(new_n631_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n439_), .A2(new_n633_), .A3(KEYINPUT43), .A4(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n632_), .A2(new_n635_), .A3(new_n595_), .A4(new_n545_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n376_), .B1(new_n637_), .B2(KEYINPUT44), .ZN(new_n638_));
  INV_X1    g437(.A(G29gat), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n636_), .B2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n529_), .B1(new_n433_), .B2(new_n440_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n545_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n596_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n585_), .A3(new_n644_), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n638_), .A2(new_n641_), .B1(new_n639_), .B2(new_n645_), .ZN(G1328gat));
  AOI21_X1  g445(.A(KEYINPUT98), .B1(new_n439_), .B2(new_n431_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n202_), .B(new_n432_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n593_), .B(new_n644_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n434_), .A2(G36gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT105), .B1(new_n649_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n642_), .A2(new_n653_), .A3(new_n644_), .A4(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n633_), .A2(KEYINPUT43), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n631_), .B(new_n658_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n439_), .A2(new_n634_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n630_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n595_), .A4(new_n545_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n636_), .A2(new_n640_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n274_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n652_), .A2(new_n654_), .A3(KEYINPUT45), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(KEYINPUT46), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n669_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n657_), .A2(new_n665_), .A3(new_n671_), .A4(new_n666_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1329gat));
  XOR2_X1   g472(.A(KEYINPUT107), .B(G43gat), .Z(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n649_), .B2(new_n352_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n662_), .A2(new_n663_), .A3(G43gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(new_n352_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g477(.A(new_n377_), .B1(new_n637_), .B2(KEYINPUT44), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n395_), .B1(new_n636_), .B2(new_n640_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n642_), .A2(new_n324_), .A3(new_n644_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n679_), .A2(new_n680_), .B1(new_n395_), .B2(new_n681_), .ZN(G1331gat));
  NOR2_X1   g481(.A1(new_n389_), .A2(new_n582_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n593_), .A2(new_n431_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G57gat), .B1(new_n686_), .B2(new_n585_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n530_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n389_), .A2(new_n431_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n598_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(KEYINPUT108), .A3(new_n598_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n376_), .A2(new_n480_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n687_), .B1(new_n695_), .B2(new_n696_), .ZN(G1332gat));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n692_), .A2(new_n274_), .A3(new_n693_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(G64gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n700_), .B1(new_n699_), .B2(G64gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n703_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(KEYINPUT48), .A3(new_n701_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n686_), .A2(new_n481_), .A3(new_n274_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n706_), .A3(new_n707_), .ZN(G1333gat));
  NAND3_X1  g507(.A1(new_n686_), .A2(new_n488_), .A3(new_n351_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G71gat), .B1(new_n694_), .B2(new_n352_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT49), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT49), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1334gat));
  INV_X1    g512(.A(KEYINPUT50), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n695_), .A2(new_n324_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G78gat), .ZN(new_n716_));
  AOI211_X1 g515(.A(KEYINPUT50), .B(new_n486_), .C1(new_n695_), .C2(new_n324_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n324_), .A2(new_n486_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT110), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n716_), .A2(new_n717_), .B1(new_n685_), .B2(new_n719_), .ZN(G1335gat));
  NAND2_X1  g519(.A1(new_n689_), .A2(new_n644_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n585_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n632_), .A2(new_n635_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n724_), .A2(KEYINPUT111), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(KEYINPUT111), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n593_), .A2(new_n431_), .A3(new_n643_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(G85gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n723_), .B1(new_n730_), .B2(new_n585_), .ZN(G1336gat));
  AOI21_X1  g530(.A(G92gat), .B1(new_n722_), .B2(new_n274_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n728_), .A2(new_n434_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n728_), .B2(new_n352_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n459_), .A2(new_n461_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n722_), .A2(new_n736_), .A3(new_n351_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT51), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n740_), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1338gat));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n632_), .A2(new_n635_), .A3(new_n324_), .A4(new_n727_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G106gat), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT52), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n748_), .A3(G106gat), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n722_), .A2(new_n444_), .A3(new_n324_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n744_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n745_), .A2(new_n748_), .A3(G106gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n748_), .B1(new_n745_), .B2(G106gat), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n744_), .B(new_n751_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n743_), .B1(new_n752_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT112), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .A3(new_n755_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n431_), .B1(new_n524_), .B2(new_n523_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n581_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n581_), .B2(new_n764_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n631_), .A2(new_n643_), .A3(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT113), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n581_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(KEYINPUT54), .A3(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n767_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  INV_X1    g572(.A(new_n495_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n491_), .A2(new_n493_), .A3(KEYINPUT66), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(KEYINPUT12), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n503_), .B1(new_n562_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n512_), .B1(new_n777_), .B2(new_n507_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n502_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n497_), .B(new_n503_), .C1(KEYINPUT12), .C2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n783_), .B2(new_n512_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(KEYINPUT114), .A3(new_n512_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n504_), .A2(KEYINPUT55), .A3(new_n505_), .A4(new_n508_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n780_), .A2(new_n784_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n519_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(KEYINPUT116), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT116), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n787_), .A2(new_n519_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT115), .B(new_n791_), .C1(new_n787_), .C2(new_n519_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n789_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n521_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n773_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n418_), .A2(KEYINPUT118), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n418_), .A2(KEYINPUT118), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n424_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n423_), .A2(new_n419_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n392_), .A3(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n430_), .A3(new_n522_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n795_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n788_), .A2(KEYINPUT116), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n793_), .A2(new_n794_), .A3(new_n792_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT117), .A3(new_n799_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n801_), .A2(new_n807_), .A3(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n596_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n596_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n793_), .A2(new_n790_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT120), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n793_), .A2(new_n819_), .A3(new_n790_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n816_), .A2(new_n818_), .A3(new_n820_), .A4(new_n821_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n806_), .A2(new_n430_), .A3(new_n521_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n822_), .A2(new_n823_), .A3(KEYINPUT58), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT58), .B1(new_n822_), .B2(new_n823_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n631_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n814_), .A2(new_n815_), .A3(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n772_), .B1(new_n827_), .B2(new_n643_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(new_n585_), .A3(new_n435_), .A4(new_n434_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n342_), .A3(new_n431_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n829_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n767_), .A2(new_n771_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n813_), .A2(new_n596_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n596_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n826_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n834_), .B1(new_n840_), .B2(new_n545_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n376_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n842_), .A2(KEYINPUT59), .A3(new_n435_), .A4(new_n434_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n432_), .B1(new_n833_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n831_), .B1(new_n844_), .B2(new_n342_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT121), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n831_), .B(new_n847_), .C1(new_n844_), .C2(new_n342_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1340gat));
  NOR3_X1   g648(.A1(new_n841_), .A2(new_n376_), .A3(new_n274_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT59), .B1(new_n850_), .B2(new_n435_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n829_), .A2(new_n832_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n530_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n833_), .A2(new_n843_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(KEYINPUT122), .A3(new_n530_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(G120gat), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n830_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(G1341gat));
  AOI21_X1  g661(.A(G127gat), .B1(new_n830_), .B2(new_n643_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n545_), .B1(new_n833_), .B2(new_n843_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g664(.A(G134gat), .B1(new_n830_), .B2(new_n597_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n856_), .A2(G134gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n634_), .ZN(G1343gat));
  NAND2_X1  g667(.A1(new_n850_), .A2(new_n436_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n432_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n688_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT123), .B(G148gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1345gat));
  NOR2_X1   g673(.A1(new_n869_), .A2(new_n545_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT61), .B(G155gat), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  INV_X1    g676(.A(G162gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n869_), .B2(new_n596_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n634_), .A2(G162gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n869_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n879_), .B(new_n883_), .C1(new_n869_), .C2(new_n880_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1347gat));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n841_), .A2(new_n585_), .A3(new_n434_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n435_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n431_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n890_), .B2(G169gat), .ZN(new_n891_));
  AOI211_X1 g690(.A(KEYINPUT62), .B(new_n222_), .C1(new_n889_), .C2(new_n431_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n432_), .A2(new_n242_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT125), .ZN(new_n894_));
  OAI22_X1  g693(.A1(new_n891_), .A2(new_n892_), .B1(new_n888_), .B2(new_n894_), .ZN(G1348gat));
  NAND3_X1  g694(.A1(new_n889_), .A2(new_n223_), .A3(new_n529_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G176gat), .B1(new_n888_), .B2(new_n688_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1349gat));
  NOR2_X1   g697(.A1(new_n888_), .A2(new_n545_), .ZN(new_n899_));
  MUX2_X1   g698(.A(G183gat), .B(new_n229_), .S(new_n899_), .Z(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n888_), .B2(new_n631_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n597_), .A2(new_n230_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n888_), .B2(new_n902_), .ZN(G1351gat));
  NAND2_X1  g702(.A1(new_n887_), .A2(new_n436_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n432_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n206_), .ZN(G1352gat));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n688_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n204_), .ZN(G1353gat));
  NOR2_X1   g707(.A1(new_n904_), .A2(new_n545_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n909_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT126), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n909_), .A2(new_n915_), .A3(new_n911_), .A4(new_n912_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT127), .B(new_n910_), .C1(new_n904_), .C2(new_n545_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n914_), .A2(new_n916_), .B1(new_n917_), .B2(new_n919_), .ZN(G1354gat));
  INV_X1    g719(.A(G218gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n904_), .A2(new_n921_), .A3(new_n631_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n887_), .A2(new_n597_), .A3(new_n436_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n921_), .B2(new_n923_), .ZN(G1355gat));
endmodule


