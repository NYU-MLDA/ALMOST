//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT31), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G71gat), .B(G99gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  OR3_X1    g008(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT82), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT81), .B(KEYINPUT26), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n216_), .A2(KEYINPUT81), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(KEYINPUT81), .ZN(new_n218_));
  OAI211_X1 g017(.A(KEYINPUT82), .B(G190gat), .C1(new_n217_), .C2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT25), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G183gat), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n215_), .A2(new_n219_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n227_), .B(KEYINPUT83), .Z(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n226_), .A2(KEYINPUT84), .A3(new_n231_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n211_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT22), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n238_), .A2(KEYINPUT85), .A3(G169gat), .ZN(new_n239_));
  INV_X1    g038(.A(G176gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(G169gat), .B1(new_n238_), .B2(KEYINPUT85), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n228_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n236_), .A2(KEYINPUT86), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT86), .ZN(new_n246_));
  INV_X1    g045(.A(new_n211_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n226_), .A2(KEYINPUT84), .A3(new_n231_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT84), .B1(new_n226_), .B2(new_n231_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n246_), .B1(new_n250_), .B2(new_n243_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT30), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n245_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT86), .B1(new_n236_), .B2(new_n244_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n246_), .A3(new_n243_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT30), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n207_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G127gat), .B(G134gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G113gat), .B(G120gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n252_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(KEYINPUT30), .A3(new_n255_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n207_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n257_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n260_), .B1(new_n257_), .B2(new_n264_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n204_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n264_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n260_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n257_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n203_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n274_));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G211gat), .B(G218gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT92), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G197gat), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n283_), .A2(G204gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(G204gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT21), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT91), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n284_), .B1(new_n287_), .B2(new_n285_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(new_n287_), .B2(new_n285_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n282_), .B(new_n286_), .C1(new_n289_), .C2(KEYINPUT21), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n281_), .A3(KEYINPUT21), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT19), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n216_), .A2(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n225_), .A2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n210_), .A2(new_n229_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT94), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(KEYINPUT94), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n227_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n298_), .B(new_n209_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT22), .B(G169gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n240_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n237_), .A2(new_n228_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT20), .B1(new_n307_), .B2(new_n292_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n294_), .A2(new_n296_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n296_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n254_), .A2(new_n293_), .A3(new_n255_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT20), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n307_), .B2(new_n292_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n310_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n279_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n296_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n292_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n308_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n310_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n278_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT100), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT100), .ZN(new_n325_));
  AOI211_X1 g124(.A(new_n325_), .B(KEYINPUT27), .C1(new_n315_), .C2(new_n321_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G155gat), .B(G162gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT89), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n328_), .A2(KEYINPUT89), .ZN(new_n330_));
  NAND3_X1  g129(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT88), .Z(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  AND2_X1   g132(.A1(KEYINPUT87), .A2(KEYINPUT2), .ZN(new_n334_));
  NOR2_X1   g133(.A1(KEYINPUT87), .A2(KEYINPUT2), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n337_));
  OR3_X1    g136(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n329_), .B(new_n330_), .C1(new_n332_), .C2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G141gat), .B(G148gat), .Z(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n341_), .B(new_n342_), .C1(KEYINPUT1), .C2(new_n328_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n292_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G233gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n347_), .A2(KEYINPUT90), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(KEYINPUT90), .ZN(new_n349_));
  OAI21_X1  g148(.A(G228gat), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n346_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n345_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G22gat), .B(G50gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT28), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n354_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n353_), .A2(new_n358_), .A3(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n344_), .A2(new_n260_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n344_), .A2(new_n260_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n365_), .ZN(new_n366_));
  OR3_X1    g165(.A1(new_n344_), .A2(KEYINPUT4), .A3(new_n260_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n363_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n376_));
  OR3_X1    g175(.A1(new_n368_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n374_), .B1(new_n368_), .B2(new_n376_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n362_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n316_), .A2(new_n296_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n310_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n279_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(KEYINPUT27), .A3(new_n321_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n327_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n378_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n366_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n364_), .A2(new_n375_), .A3(new_n365_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n373_), .A3(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n378_), .B2(new_n386_), .ZN(new_n391_));
  OR3_X1    g190(.A1(new_n322_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(KEYINPUT32), .B(new_n278_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT99), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n278_), .A2(KEYINPUT32), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT98), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n317_), .A2(new_n320_), .A3(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n393_), .A2(new_n379_), .A3(new_n394_), .A4(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n379_), .A3(new_n397_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT99), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n392_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n362_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n273_), .B1(new_n385_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n384_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT101), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT101), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n384_), .B(new_n406_), .C1(new_n324_), .C2(new_n326_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n379_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n273_), .A2(new_n408_), .A3(new_n362_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT102), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT102), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n405_), .A2(new_n409_), .A3(new_n412_), .A4(new_n407_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n403_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G43gat), .B(G50gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT72), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(G29gat), .ZN(new_n417_));
  INV_X1    g216(.A(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT15), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n417_), .B(G36gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT15), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT64), .B(G92gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G85gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n425_), .A2(new_n426_), .B1(KEYINPUT9), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G99gat), .A2(G106gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT6), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT10), .B(G99gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(G106gat), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n433_), .B(KEYINPUT65), .Z(new_n434_));
  INV_X1    g233(.A(KEYINPUT8), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n436_));
  INV_X1    g235(.A(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G106gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n429_), .B(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n443_), .B2(KEYINPUT68), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(KEYINPUT68), .B2(new_n443_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n427_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n435_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n430_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n449_), .A2(KEYINPUT66), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(KEYINPUT66), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n435_), .B(new_n447_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n452_), .B2(KEYINPUT67), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n435_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(KEYINPUT66), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n453_), .A2(new_n459_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n420_), .A2(new_n423_), .B1(new_n434_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G232gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT71), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT34), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT35), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n460_), .A2(new_n434_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(new_n421_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n465_), .A2(new_n466_), .ZN(new_n470_));
  OR3_X1    g269(.A1(new_n461_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G190gat), .B(G218gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G134gat), .B(G162gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(KEYINPUT36), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n470_), .B1(new_n461_), .B2(new_n469_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n471_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n474_), .B(KEYINPUT36), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT105), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n414_), .A2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n483_), .A2(KEYINPUT106), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(KEYINPUT106), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G230gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G71gat), .B(G78gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(G57gat), .B(G64gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(KEYINPUT11), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(KEYINPUT11), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n468_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n445_), .A2(new_n447_), .ZN(new_n496_));
  OAI22_X1  g295(.A1(new_n457_), .A2(new_n458_), .B1(new_n496_), .B2(new_n435_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n452_), .A2(KEYINPUT67), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n434_), .B(new_n495_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(KEYINPUT12), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(KEYINPUT12), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n495_), .B1(new_n460_), .B2(new_n434_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n488_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n487_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT70), .ZN(new_n507_));
  XOR2_X1   g306(.A(G120gat), .B(G148gat), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G176gat), .B(G204gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  OR3_X1    g310(.A1(new_n504_), .A2(new_n505_), .A3(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n515_), .A2(KEYINPUT13), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(KEYINPUT13), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT75), .B(G15gat), .ZN(new_n520_));
  INV_X1    g319(.A(G22gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(G1gat), .ZN(new_n523_));
  INV_X1    g322(.A(G8gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G8gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT76), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(new_n495_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G183gat), .B(G211gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G127gat), .B(G155gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT17), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n532_), .A2(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n539_), .A2(KEYINPUT78), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(KEYINPUT78), .A3(new_n538_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n532_), .A2(new_n542_), .A3(new_n537_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n540_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n420_), .A2(new_n423_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n528_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n421_), .A2(new_n528_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n421_), .B(new_n528_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n546_), .A2(new_n550_), .B1(new_n551_), .B2(new_n549_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(G169gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n283_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT80), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT80), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n552_), .A2(new_n558_), .A3(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n552_), .A2(new_n555_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n519_), .A2(new_n544_), .A3(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n486_), .A2(new_n379_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(G1gat), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n477_), .A2(KEYINPUT73), .B1(new_n480_), .B2(KEYINPUT74), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n480_), .A2(KEYINPUT74), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT37), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n480_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n471_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n571_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n544_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n518_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT79), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n414_), .A2(new_n563_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n581_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT103), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT103), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n582_), .A2(new_n583_), .A3(new_n587_), .A4(new_n584_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n586_), .A2(new_n523_), .A3(new_n379_), .A4(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n589_), .A2(KEYINPUT104), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(KEYINPUT104), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n566_), .B1(new_n593_), .B2(new_n594_), .ZN(G1324gat));
  AND2_X1   g394(.A1(new_n586_), .A2(new_n588_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n405_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n407_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(new_n524_), .A3(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n600_), .B(new_n564_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n602_), .A2(new_n603_), .A3(G8gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n602_), .B2(G8gat), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n601_), .B(KEYINPUT40), .C1(new_n604_), .C2(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1325gat));
  INV_X1    g409(.A(G15gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n596_), .A2(new_n611_), .A3(new_n273_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n486_), .A2(new_n273_), .A3(new_n564_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n613_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT41), .B1(new_n613_), .B2(G15gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(G1326gat));
  INV_X1    g415(.A(new_n362_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n596_), .A2(new_n521_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n486_), .A2(new_n617_), .A3(new_n564_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G22gat), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(KEYINPUT42), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(KEYINPUT42), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n618_), .B1(new_n621_), .B2(new_n622_), .ZN(G1327gat));
  NAND2_X1  g422(.A1(new_n482_), .A2(new_n544_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT109), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n519_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n583_), .ZN(new_n627_));
  INV_X1    g426(.A(G29gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n379_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n519_), .A2(new_n579_), .A3(new_n563_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n411_), .A2(new_n413_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n403_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT107), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n570_), .A2(new_n635_), .A3(new_n577_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n571_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT107), .B1(new_n637_), .B2(new_n576_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n631_), .B1(new_n634_), .B2(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n414_), .A2(KEYINPUT43), .A3(new_n578_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n630_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n630_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n578_), .A2(KEYINPUT43), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n634_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT43), .B1(new_n414_), .B2(new_n639_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT44), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n379_), .A3(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT108), .B1(new_n652_), .B2(G29gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n629_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  NAND4_X1  g455(.A1(new_n626_), .A2(new_n418_), .A3(new_n600_), .A4(new_n583_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT45), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n645_), .A2(new_n600_), .A3(new_n651_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(new_n418_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n658_), .B(KEYINPUT46), .C1(new_n418_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  AND2_X1   g463(.A1(new_n627_), .A2(new_n273_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n645_), .A2(G43gat), .A3(new_n273_), .ZN(new_n666_));
  AOI211_X1 g465(.A(new_n644_), .B(new_n646_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n667_));
  OAI22_X1  g466(.A1(G43gat), .A2(new_n665_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g468(.A(KEYINPUT110), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n617_), .B1(new_n650_), .B2(KEYINPUT44), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n667_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n645_), .A2(KEYINPUT110), .A3(new_n651_), .A4(new_n617_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(G50gat), .ZN(new_n674_));
  INV_X1    g473(.A(G50gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n627_), .A2(new_n675_), .A3(new_n617_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT111), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n674_), .A2(KEYINPUT111), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1331gat));
  NOR2_X1   g480(.A1(new_n518_), .A2(new_n562_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n634_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n637_), .A2(new_n576_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(new_n544_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n379_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT112), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n518_), .A2(new_n544_), .A3(new_n562_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n486_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n379_), .A2(G57gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1332gat));
  INV_X1    g491(.A(G64gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n685_), .A2(new_n693_), .A3(new_n600_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G64gat), .B1(new_n689_), .B2(new_n599_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT48), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT48), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(G1333gat));
  INV_X1    g497(.A(new_n273_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(G71gat), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT113), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n685_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G71gat), .B1(new_n689_), .B2(new_n699_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT49), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT49), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(G1334gat));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n685_), .A2(new_n707_), .A3(new_n617_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G78gat), .B1(new_n689_), .B2(new_n362_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(G1335gat));
  NOR2_X1   g511(.A1(new_n683_), .A2(new_n625_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n379_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n682_), .A2(new_n544_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT114), .Z(new_n717_));
  AND2_X1   g516(.A1(new_n379_), .A2(G85gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1336gat));
  AOI21_X1  g518(.A(G92gat), .B1(new_n713_), .B2(new_n600_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n600_), .A2(new_n424_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n717_), .B2(new_n721_), .ZN(G1337gat));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n273_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G99gat), .ZN(new_n724_));
  INV_X1    g523(.A(new_n431_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n713_), .A2(new_n725_), .A3(new_n273_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727_));
  AOI22_X1  g526(.A1(new_n724_), .A2(new_n726_), .B1(KEYINPUT115), .B2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(KEYINPUT115), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(G1338gat));
  INV_X1    g529(.A(KEYINPUT116), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  OAI21_X1  g531(.A(G106gat), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n716_), .B2(new_n617_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n732_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n713_), .A2(new_n438_), .A3(new_n617_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1339gat));
  NAND4_X1  g540(.A1(new_n578_), .A2(new_n518_), .A3(new_n579_), .A4(new_n563_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n482_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n562_), .A2(new_n512_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n511_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n500_), .A2(new_n503_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT55), .B1(new_n748_), .B2(new_n487_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n750_), .B(new_n488_), .C1(new_n500_), .C2(new_n503_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n500_), .A2(new_n488_), .A3(new_n503_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n500_), .A2(new_n503_), .A3(KEYINPUT117), .A4(new_n488_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n747_), .B1(new_n752_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT118), .B1(new_n758_), .B2(KEYINPUT56), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n755_), .A2(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n504_), .A2(KEYINPUT55), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n501_), .A2(new_n502_), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT12), .B(new_n495_), .C1(new_n460_), .C2(new_n434_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n487_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n750_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n761_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n511_), .B1(new_n760_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n759_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT119), .B1(new_n758_), .B2(KEYINPUT56), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n757_), .A2(new_n765_), .A3(new_n761_), .ZN(new_n773_));
  AND4_X1   g572(.A1(KEYINPUT119), .A2(new_n773_), .A3(KEYINPUT56), .A4(new_n511_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n746_), .B1(new_n771_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n551_), .A2(new_n548_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n555_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(KEYINPUT120), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT120), .B1(new_n777_), .B2(new_n778_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n547_), .A2(new_n548_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n546_), .B2(new_n781_), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n779_), .A2(new_n782_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n514_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT57), .B(new_n745_), .C1(new_n776_), .C2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n511_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n758_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n759_), .A2(new_n789_), .A3(new_n770_), .A4(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n746_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n784_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n786_), .B1(new_n793_), .B2(new_n482_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n783_), .A2(new_n512_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n767_), .A2(new_n769_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n787_), .B2(new_n796_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n797_), .A2(KEYINPUT58), .ZN(new_n798_));
  INV_X1    g597(.A(new_n795_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n787_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n758_), .A2(KEYINPUT56), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n799_), .B(KEYINPUT58), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n798_), .A2(new_n684_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n785_), .A2(new_n794_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n744_), .B1(new_n804_), .B2(new_n544_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n699_), .A2(new_n617_), .A3(new_n408_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n599_), .A2(new_n806_), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n805_), .A2(KEYINPUT59), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT121), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n798_), .A2(new_n809_), .A3(new_n684_), .A4(new_n802_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n684_), .B1(new_n797_), .B2(KEYINPUT58), .ZN(new_n811_));
  INV_X1    g610(.A(new_n802_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT121), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n785_), .A2(new_n794_), .A3(new_n810_), .A4(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n744_), .B1(new_n814_), .B2(new_n544_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT59), .B1(new_n815_), .B2(new_n807_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n817_));
  INV_X1    g616(.A(G113gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n563_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n808_), .A2(new_n816_), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(G113gat), .B1(new_n820_), .B2(KEYINPUT122), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n815_), .A2(new_n807_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n562_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1340gat));
  NAND2_X1  g623(.A1(new_n814_), .A2(new_n544_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n744_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n807_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n518_), .A2(G120gat), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n827_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n519_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n808_), .A2(new_n816_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G120gat), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n830_), .A2(KEYINPUT60), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1341gat));
  OAI21_X1  g634(.A(G127gat), .B1(new_n832_), .B2(new_n544_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n822_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n544_), .A2(G127gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1342gat));
  OAI21_X1  g638(.A(G134gat), .B1(new_n832_), .B2(new_n578_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n745_), .A2(G134gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n837_), .B2(new_n841_), .ZN(G1343gat));
  NOR4_X1   g641(.A1(new_n600_), .A2(new_n408_), .A3(new_n362_), .A4(new_n273_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n827_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n562_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT123), .B(G141gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1344gat));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n519_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g649(.A1(new_n845_), .A2(new_n579_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  AND3_X1   g652(.A1(new_n845_), .A2(G162gat), .A3(new_n640_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G162gat), .B1(new_n845_), .B2(new_n482_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1347gat));
  INV_X1    g655(.A(new_n409_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n599_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n805_), .A2(new_n563_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G169gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n863_));
  OR3_X1    g662(.A1(new_n860_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n304_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(G1348gat));
  NOR2_X1   g666(.A1(new_n518_), .A2(new_n240_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n815_), .A2(new_n859_), .A3(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n805_), .A2(new_n518_), .A3(new_n859_), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n870_), .A2(KEYINPUT125), .B1(new_n871_), .B2(G176gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n827_), .A2(new_n858_), .A3(new_n868_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT126), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n871_), .A2(G176gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n870_), .A2(KEYINPUT125), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n877_), .A2(new_n878_), .A3(new_n879_), .A4(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n881_), .ZN(G1349gat));
  NAND3_X1  g681(.A1(new_n827_), .A2(new_n579_), .A3(new_n858_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n805_), .A2(new_n859_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n544_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n883_), .A2(new_n221_), .B1(new_n884_), .B2(new_n885_), .ZN(G1350gat));
  NAND4_X1  g685(.A1(new_n884_), .A2(new_n482_), .A3(new_n220_), .A4(new_n297_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n805_), .A2(new_n578_), .A3(new_n859_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n214_), .ZN(G1351gat));
  NOR4_X1   g688(.A1(new_n599_), .A2(new_n379_), .A3(new_n362_), .A4(new_n273_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n827_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n563_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n283_), .ZN(G1352gat));
  INV_X1    g692(.A(new_n891_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n519_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT127), .B(G204gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1353gat));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  AND2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n891_), .A2(new_n544_), .A3(new_n898_), .A4(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n894_), .A2(new_n579_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n898_), .ZN(G1354gat));
  OR3_X1    g701(.A1(new_n891_), .A2(G218gat), .A3(new_n745_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G218gat), .B1(new_n891_), .B2(new_n578_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1355gat));
endmodule


