//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G231gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G57gat), .B(G64gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT11), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(KEYINPUT11), .ZN(new_n213_));
  XOR2_X1   g012(.A(G71gat), .B(G78gat), .Z(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n210_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT16), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(G211gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G127gat), .B(G155gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n219_), .B(new_n220_), .Z(new_n221_));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n217_), .B1(KEYINPUT70), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n221_), .B(KEYINPUT17), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT78), .ZN(new_n227_));
  INV_X1    g026(.A(new_n223_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n217_), .B1(KEYINPUT70), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n225_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT73), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G29gat), .B(G36gat), .ZN(new_n233_));
  INV_X1    g032(.A(G43gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G50gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n233_), .B(G43gat), .ZN(new_n237_));
  INV_X1    g036(.A(G50gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT15), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT15), .B1(new_n236_), .B2(new_n239_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT10), .B(G99gat), .Z(new_n245_));
  INV_X1    g044(.A(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT65), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G99gat), .A2(G106gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT6), .ZN(new_n250_));
  INV_X1    g049(.A(G85gat), .ZN(new_n251_));
  INV_X1    g050(.A(G92gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT9), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G85gat), .B(G92gat), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT9), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n245_), .A2(new_n259_), .A3(new_n246_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n248_), .A2(new_n256_), .A3(new_n258_), .A4(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n258_), .A2(new_n250_), .A3(new_n255_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(KEYINPUT69), .A3(new_n248_), .A4(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n257_), .A2(KEYINPUT67), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G85gat), .A2(G92gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n253_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n272_));
  OR3_X1    g071(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n250_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n272_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT8), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT66), .B1(new_n267_), .B2(new_n270_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT8), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n275_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n266_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n232_), .B1(new_n244_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n242_), .A2(new_n243_), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n263_), .A2(new_n265_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n284_), .A2(new_n285_), .A3(KEYINPUT73), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT74), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n248_), .A2(new_n260_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n277_), .A2(new_n280_), .B1(new_n264_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n244_), .A2(new_n232_), .A3(new_n282_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT73), .B1(new_n284_), .B2(new_n285_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n287_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT34), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n297_), .A2(KEYINPUT35), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G190gat), .B(G218gat), .ZN(new_n300_));
  INV_X1    g099(.A(G134gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G162gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT36), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n297_), .A2(KEYINPUT35), .ZN(new_n306_));
  AOI211_X1 g105(.A(new_n298_), .B(new_n306_), .C1(new_n291_), .C2(new_n293_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n290_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n299_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n303_), .B(new_n304_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n295_), .A2(new_n298_), .B1(new_n290_), .B2(new_n307_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n309_), .B(new_n310_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT37), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT37), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT75), .B1(new_n312_), .B2(new_n311_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n316_), .A2(KEYINPUT75), .B1(new_n317_), .B2(new_n309_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT77), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n313_), .A2(new_n314_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n316_), .A2(KEYINPUT75), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n317_), .A2(new_n309_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n320_), .B(new_n321_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n231_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n216_), .B(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n282_), .A2(KEYINPUT12), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G230gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT64), .ZN(new_n330_));
  INV_X1    g129(.A(new_n280_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n279_), .B1(new_n278_), .B2(new_n275_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n261_), .B(new_n216_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT12), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n289_), .B2(new_n216_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n328_), .A2(new_n330_), .A3(new_n333_), .A4(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n289_), .A2(KEYINPUT68), .A3(new_n216_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n289_), .A2(new_n216_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n330_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G120gat), .B(G148gat), .ZN(new_n344_));
  INV_X1    g143(.A(G204gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT5), .ZN(new_n347_));
  INV_X1    g146(.A(G176gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n337_), .A2(new_n343_), .A3(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n350_), .B1(new_n337_), .B2(new_n343_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT13), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n325_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT79), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n206_), .B(new_n207_), .Z(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n240_), .A2(new_n208_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(G229gat), .A3(G233gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n244_), .A2(new_n208_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G229gat), .A2(G233gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n368_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G113gat), .B(G141gat), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G197gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n373_), .A2(new_n376_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n366_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(KEYINPUT81), .A3(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G15gat), .B(G43gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT86), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n393_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G183gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT82), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G183gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT25), .ZN(new_n401_));
  OR2_X1    g200(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G190gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT26), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT83), .B1(new_n404_), .B2(KEYINPUT26), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT26), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(G190gat), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n403_), .A2(new_n405_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT84), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n378_), .A2(new_n348_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT24), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G169gat), .A2(G176gat), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G183gat), .A2(G190gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT23), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT85), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n417_), .A2(new_n420_), .A3(new_n424_), .A4(new_n421_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n416_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n405_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n410_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n412_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n420_), .A2(new_n421_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n398_), .A2(new_n400_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(G190gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT22), .B(G169gat), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n413_), .B1(new_n436_), .B2(new_n348_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n431_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT30), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n440_), .A2(new_n441_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n396_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n442_), .B2(new_n396_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G127gat), .A2(G134gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G127gat), .A2(G134gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(G113gat), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(G127gat), .A2(G134gat), .ZN(new_n450_));
  INV_X1    g249(.A(G113gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G120gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(G120gat), .B1(new_n449_), .B2(new_n452_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT31), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n445_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n445_), .A2(new_n459_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n453_), .B(new_n454_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G155gat), .B(G162gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT3), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT2), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT88), .B1(G141gat), .B2(G148gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n470_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n474_), .A2(new_n475_), .A3(new_n472_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n465_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n465_), .A2(KEYINPUT1), .ZN(new_n480_));
  INV_X1    g279(.A(new_n466_), .ZN(new_n481_));
  AND2_X1   g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n482_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n464_), .B1(new_n479_), .B2(new_n485_), .ZN(new_n486_));
  OAI22_X1  g285(.A1(new_n475_), .A2(new_n474_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n478_), .A2(new_n487_), .A3(new_n469_), .A4(new_n468_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n465_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n457_), .A2(new_n490_), .A3(new_n484_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n486_), .A2(new_n491_), .A3(KEYINPUT4), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G225gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n484_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT4), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n464_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n486_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G1gat), .B(G29gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(G57gat), .B(G85gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(new_n505_), .A3(new_n499_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT18), .B(G64gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(G92gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G8gat), .B(G36gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n380_), .A2(G204gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n345_), .B2(G197gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n380_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n515_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT21), .ZN(new_n522_));
  XOR2_X1   g321(.A(G211gat), .B(G218gat), .Z(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT25), .B(G183gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G190gat), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n416_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n422_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n433_), .B1(G183gat), .B2(G190gat), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n528_), .A2(new_n529_), .B1(new_n530_), .B2(new_n437_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G197gat), .B(G204gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT21), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT90), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n345_), .A2(G197gat), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n535_), .B(KEYINPUT21), .C1(new_n515_), .C2(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n523_), .B1(new_n519_), .B2(new_n533_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT92), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n515_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n380_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT91), .B1(new_n380_), .B2(G204gat), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n541_), .B(new_n533_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n523_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(new_n534_), .A3(new_n545_), .A4(new_n537_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n525_), .B(new_n531_), .C1(new_n540_), .C2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n438_), .ZN(new_n550_));
  AND4_X1   g349(.A1(new_n429_), .A2(new_n403_), .A3(new_n405_), .A4(new_n410_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n429_), .B1(new_n428_), .B2(new_n410_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n553_), .B2(new_n426_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n522_), .A2(new_n524_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n538_), .A2(KEYINPUT92), .A3(new_n539_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n546_), .A2(new_n547_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n555_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n549_), .B(KEYINPUT20), .C1(new_n554_), .C2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G226gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT19), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT20), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n525_), .B1(new_n540_), .B2(new_n548_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n531_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n554_), .A2(new_n558_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n563_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n514_), .B1(new_n562_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT20), .B1(new_n558_), .B2(new_n531_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n565_), .A2(new_n439_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n561_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n564_), .B1(new_n565_), .B2(new_n439_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n563_), .A3(new_n549_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n514_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n570_), .A2(new_n571_), .A3(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n574_), .A2(new_n576_), .A3(KEYINPUT95), .A4(new_n577_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT27), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n572_), .A2(new_n573_), .A3(new_n561_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n563_), .B1(new_n575_), .B2(new_n549_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n514_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(KEYINPUT27), .A3(new_n578_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n495_), .A2(KEYINPUT29), .ZN(new_n588_));
  OAI211_X1 g387(.A(G228gat), .B(G233gat), .C1(new_n588_), .C2(new_n558_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G228gat), .A2(G233gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n495_), .A2(KEYINPUT29), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n565_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G78gat), .B(G106gat), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n495_), .A2(KEYINPUT29), .ZN(new_n597_));
  XOR2_X1   g396(.A(G22gat), .B(G50gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT28), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n597_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n589_), .A2(new_n592_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n593_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n594_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n601_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n587_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n463_), .A2(new_n510_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n577_), .A2(KEYINPUT32), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n574_), .A2(new_n576_), .A3(new_n610_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n509_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n579_), .A2(new_n580_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n508_), .A2(KEYINPUT33), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n498_), .A2(new_n617_), .A3(new_n505_), .A4(new_n499_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n486_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n491_), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n620_), .A2(new_n621_), .A3(KEYINPUT97), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT97), .B1(new_n620_), .B2(new_n621_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n494_), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n492_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n506_), .A3(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n619_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n614_), .B1(new_n615_), .B2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT98), .B1(new_n628_), .B2(new_n606_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n606_), .A2(new_n510_), .A3(new_n582_), .A4(new_n586_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n601_), .A2(new_n605_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n601_), .A2(new_n605_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n619_), .A2(new_n626_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n580_), .B2(new_n579_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n633_), .B(new_n634_), .C1(new_n636_), .C2(new_n614_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n629_), .A2(new_n630_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n462_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(KEYINPUT99), .A3(new_n462_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n609_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n365_), .A2(new_n390_), .A3(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n509_), .B(KEYINPUT100), .Z(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n203_), .A3(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT38), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n638_), .A2(KEYINPUT99), .A3(new_n462_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT99), .B1(new_n638_), .B2(new_n462_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n608_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n362_), .A2(new_n390_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n309_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n231_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n510_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n648_), .A2(new_n659_), .ZN(G1324gat));
  AOI21_X1  g459(.A(new_n204_), .B1(new_n657_), .B2(new_n587_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT39), .Z(new_n662_));
  NAND3_X1  g461(.A1(new_n644_), .A2(new_n204_), .A3(new_n587_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n662_), .A2(KEYINPUT40), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n657_), .B2(new_n463_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT41), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n644_), .A2(new_n669_), .A3(new_n463_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1326gat));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n657_), .B2(new_n606_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT42), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n644_), .A2(new_n674_), .A3(new_n606_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n319_), .A2(new_n324_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n651_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n651_), .B2(new_n680_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n231_), .B(new_n652_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n319_), .A2(new_n324_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n643_), .B2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n651_), .A2(new_n680_), .A3(new_n679_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n689_), .A2(KEYINPUT44), .A3(new_n231_), .A4(new_n652_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n685_), .A2(new_n646_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G29gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n654_), .A2(new_n230_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT101), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n653_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n510_), .A2(G29gat), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT102), .Z(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n692_), .A2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n695_), .A2(new_n700_), .A3(new_n701_), .A4(new_n587_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n653_), .A2(new_n701_), .A3(new_n694_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n587_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT103), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n702_), .A2(KEYINPUT45), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT45), .B1(new_n702_), .B2(new_n705_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n685_), .A2(new_n587_), .A3(new_n690_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n708_), .B(new_n710_), .C1(KEYINPUT104), .C2(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1329gat));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n685_), .A2(G43gat), .A3(new_n463_), .A4(new_n690_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n695_), .A2(new_n463_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n234_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n718_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n718_), .B1(new_n717_), .B2(new_n720_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n716_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n723_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(KEYINPUT47), .A3(new_n721_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  NAND3_X1  g526(.A1(new_n695_), .A2(new_n238_), .A3(new_n606_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n685_), .A2(new_n606_), .A3(new_n690_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n729_), .A2(KEYINPUT106), .A3(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT106), .B1(new_n729_), .B2(G50gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(G1331gat));
  NAND2_X1  g531(.A1(new_n325_), .A2(new_n362_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n733_), .A2(KEYINPUT107), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(KEYINPUT107), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n641_), .A2(new_n642_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n389_), .B1(new_n736_), .B2(new_n608_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(new_n645_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(G57gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n656_), .A3(new_n362_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(new_n510_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(G57gat), .B2(new_n742_), .ZN(G1332gat));
  OAI21_X1  g542(.A(G64gat), .B1(new_n741_), .B2(new_n704_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT48), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n704_), .A2(G64gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n738_), .B2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n741_), .B2(new_n462_), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT109), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n748_), .B(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n462_), .A2(G71gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n738_), .B2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n741_), .B2(new_n633_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n633_), .A2(G78gat), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT110), .Z(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n738_), .B2(new_n757_), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n389_), .A2(new_n230_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n362_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n762_), .A2(new_n251_), .A3(new_n510_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n737_), .A2(new_n764_), .A3(new_n362_), .A4(new_n694_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n651_), .A2(new_n390_), .A3(new_n362_), .A4(new_n694_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT111), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n646_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n763_), .A2(new_n769_), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n762_), .A2(new_n252_), .A3(new_n704_), .ZN(new_n771_));
  AOI21_X1  g570(.A(G92gat), .B1(new_n768_), .B2(new_n587_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1337gat));
  INV_X1    g572(.A(new_n760_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n463_), .B(new_n774_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G99gat), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n463_), .A2(new_n245_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n766_), .A2(KEYINPUT111), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n766_), .A2(KEYINPUT111), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n776_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT112), .B1(new_n782_), .B2(KEYINPUT51), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n784_), .B(new_n785_), .C1(new_n776_), .C2(new_n781_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n768_), .A2(new_n778_), .B1(new_n775_), .B2(G99gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT113), .B1(new_n787_), .B2(new_n785_), .ZN(new_n788_));
  INV_X1    g587(.A(G99gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n761_), .B2(new_n463_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n777_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  NOR4_X1   g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .A4(KEYINPUT51), .ZN(new_n793_));
  OAI22_X1  g592(.A1(new_n783_), .A2(new_n786_), .B1(new_n788_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n784_), .B1(new_n787_), .B2(new_n785_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n782_), .A2(KEYINPUT112), .A3(KEYINPUT51), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(KEYINPUT114), .C1(new_n788_), .C2(new_n793_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n796_), .A2(new_n800_), .ZN(G1338gat));
  NAND3_X1  g600(.A1(new_n768_), .A2(new_n246_), .A3(new_n606_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n761_), .A2(new_n606_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G106gat), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n336_), .B2(KEYINPUT116), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n336_), .B2(new_n809_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n341_), .A2(new_n335_), .A3(new_n328_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n341_), .A2(KEYINPUT117), .A3(new_n335_), .A4(new_n328_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n330_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n809_), .B(new_n811_), .C1(new_n336_), .C2(KEYINPUT116), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n813_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n349_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n810_), .A2(new_n812_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n816_), .A2(new_n817_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n330_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n819_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n822_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n350_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n821_), .A2(new_n351_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  AND4_X1   g630(.A1(G229gat), .A2(new_n374_), .A3(G233gat), .A4(new_n368_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n375_), .B2(new_n372_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n384_), .B1(new_n833_), .B2(new_n381_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n830_), .A2(new_n831_), .A3(KEYINPUT58), .A4(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n821_), .A2(new_n829_), .A3(new_n351_), .A4(new_n834_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT120), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n837_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n319_), .A2(new_n324_), .A3(new_n840_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n821_), .A2(new_n829_), .A3(new_n389_), .A4(new_n351_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n834_), .A2(new_n353_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n654_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n845_), .A2(KEYINPUT119), .A3(new_n654_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n845_), .A2(KEYINPUT57), .A3(new_n654_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n842_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n231_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n390_), .B(new_n230_), .C1(new_n357_), .C2(new_n359_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT115), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n686_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n686_), .B2(new_n856_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n854_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n463_), .A2(new_n607_), .A3(new_n646_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866_), .B2(new_n389_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT119), .B1(new_n845_), .B2(new_n654_), .ZN(new_n868_));
  AOI211_X1 g667(.A(new_n847_), .B(new_n655_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n868_), .A2(new_n869_), .A3(KEYINPUT57), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n839_), .A2(new_n841_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT121), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n842_), .A2(new_n851_), .A3(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n874_), .A3(new_n852_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n231_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n861_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n863_), .A2(KEYINPUT59), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n877_), .A2(new_n878_), .B1(new_n865_), .B2(KEYINPUT59), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n389_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n867_), .B1(new_n881_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g681(.A(new_n454_), .B1(new_n363_), .B2(KEYINPUT60), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n866_), .B(new_n883_), .C1(KEYINPUT60), .C2(new_n454_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n362_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n886_), .B2(new_n454_), .ZN(G1341gat));
  AOI21_X1  g686(.A(G127gat), .B1(new_n866_), .B2(new_n230_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n230_), .A2(G127gat), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT122), .Z(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n879_), .B2(new_n890_), .ZN(G1342gat));
  OAI21_X1  g690(.A(new_n301_), .B1(new_n865_), .B2(new_n654_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n860_), .B1(new_n853_), .B2(new_n231_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT59), .B1(new_n893_), .B2(new_n863_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n860_), .B1(new_n875_), .B2(new_n231_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n878_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n894_), .B(G134gat), .C1(new_n895_), .C2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n892_), .B1(new_n897_), .B2(new_n686_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT123), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n900_), .B(new_n892_), .C1(new_n897_), .C2(new_n686_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1343gat));
  NOR3_X1   g701(.A1(new_n893_), .A2(new_n463_), .A3(new_n645_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n587_), .A2(new_n633_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n389_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n362_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n230_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT61), .B(G155gat), .Z(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT124), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n910_), .B(new_n912_), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n905_), .B2(new_n655_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n680_), .A2(G162gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT125), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n905_), .B2(new_n916_), .ZN(G1347gat));
  NOR3_X1   g716(.A1(new_n462_), .A2(new_n704_), .A3(new_n646_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n877_), .A2(new_n389_), .A3(new_n633_), .A4(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n919_), .A2(new_n920_), .A3(G169gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n919_), .B2(G169gat), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n895_), .A2(new_n606_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n918_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n389_), .A2(new_n436_), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT126), .Z(new_n926_));
  OAI22_X1  g725(.A1(new_n921_), .A2(new_n922_), .B1(new_n924_), .B2(new_n926_), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n923_), .A2(new_n362_), .A3(new_n918_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n893_), .A2(new_n606_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n918_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n363_), .A2(new_n348_), .A3(new_n930_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n928_), .A2(new_n348_), .B1(new_n929_), .B2(new_n931_), .ZN(G1349gat));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n231_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n434_), .B1(new_n929_), .B2(new_n933_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n930_), .A2(new_n231_), .A3(new_n526_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n923_), .B2(new_n935_), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n924_), .B2(new_n686_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n655_), .A2(new_n527_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n924_), .B2(new_n938_), .ZN(G1351gat));
  NOR2_X1   g738(.A1(new_n633_), .A2(new_n509_), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n862_), .A2(new_n462_), .A3(new_n940_), .A4(new_n587_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n390_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n380_), .ZN(G1352gat));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n363_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(new_n345_), .ZN(G1353gat));
  NOR2_X1   g744(.A1(new_n941_), .A2(new_n231_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n946_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT63), .B(G211gat), .Z(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n946_), .B2(new_n948_), .ZN(G1354gat));
  INV_X1    g748(.A(G218gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n941_), .A2(new_n950_), .A3(new_n686_), .ZN(new_n951_));
  NOR4_X1   g750(.A1(new_n893_), .A2(new_n509_), .A3(new_n463_), .A4(new_n633_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n952_), .A2(new_n953_), .A3(new_n655_), .A4(new_n587_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT127), .B1(new_n941_), .B2(new_n654_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n951_), .B1(new_n956_), .B2(new_n950_), .ZN(G1355gat));
endmodule


