//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  OR3_X1    g001(.A1(new_n202_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT87), .B1(new_n202_), .B2(KEYINPUT1), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .A4(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n205_), .A2(new_n202_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT88), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n210_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT88), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n209_), .A2(new_n216_), .B1(new_n217_), .B2(KEYINPUT3), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(new_n216_), .B2(new_n209_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n212_), .B1(new_n215_), .B2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n220_), .A2(KEYINPUT89), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(KEYINPUT89), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n211_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n220_), .B(KEYINPUT89), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(new_n226_), .A3(new_n211_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G225gat), .A2(G233gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n228_), .A2(KEYINPUT4), .A3(new_n230_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n232_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n223_), .A2(new_n236_), .A3(new_n227_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G1gat), .B(G29gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G85gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G57gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n233_), .A2(new_n238_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT86), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G71gat), .B(G99gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(G43gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n251_), .B(new_n253_), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT23), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(G183gat), .A3(G190gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G183gat), .ZN(new_n260_));
  INV_X1    g059(.A(G190gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT23), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n258_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT25), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(G183gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT25), .B(G183gat), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT82), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT24), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n265_), .B1(new_n279_), .B2(KEYINPUT83), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n276_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n277_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT83), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n262_), .A2(new_n257_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(G183gat), .B2(G190gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(KEYINPUT22), .B(G169gat), .Z(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(G176gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(new_n274_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n280_), .A2(new_n285_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n287_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n281_), .B1(new_n279_), .B2(KEYINPUT83), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n264_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(KEYINPUT30), .ZN(new_n298_));
  OAI21_X1  g097(.A(G15gat), .B1(new_n293_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n291_), .A2(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(KEYINPUT30), .ZN(new_n301_));
  INV_X1    g100(.A(G15gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n299_), .A2(new_n227_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n227_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n255_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n226_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n299_), .A2(new_n227_), .A3(new_n303_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n254_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G78gat), .B(G106gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n223_), .A2(KEYINPUT29), .ZN(new_n313_));
  XOR2_X1   g112(.A(G211gat), .B(G218gat), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT91), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT91), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G197gat), .B(G204gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT92), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT21), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n321_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n319_), .A2(KEYINPUT93), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT93), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n315_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(new_n322_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n319_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT90), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n320_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT21), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G228gat), .ZN(new_n337_));
  INV_X1    g136(.A(G233gat), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n313_), .B(new_n336_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n338_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n229_), .B2(new_n211_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n325_), .A2(new_n328_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n340_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G22gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n339_), .B2(new_n344_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n312_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n339_), .A2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G22gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n312_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n346_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n229_), .A2(new_n341_), .A3(new_n211_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n354_), .A2(KEYINPUT28), .ZN(new_n355_));
  INV_X1    g154(.A(G50gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(KEYINPUT28), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n349_), .A2(new_n353_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n311_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n349_), .A2(new_n353_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n360_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n306_), .A2(new_n310_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n349_), .A2(new_n353_), .A3(new_n360_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n247_), .B1(new_n363_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT94), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n291_), .A2(new_n343_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(KEYINPUT20), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  AOI211_X1 g174(.A(KEYINPUT94), .B(new_n375_), .C1(new_n291_), .C2(new_n343_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT101), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT19), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n382_));
  INV_X1    g181(.A(new_n286_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n383_), .B2(new_n282_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n271_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n266_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n286_), .A2(KEYINPUT95), .A3(new_n281_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n384_), .A2(new_n278_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n290_), .B1(new_n265_), .B2(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n390_), .A2(KEYINPUT96), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(KEYINPUT96), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n336_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n377_), .A2(new_n378_), .A3(new_n381_), .A4(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n297_), .B2(new_n336_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT94), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n373_), .A2(new_n372_), .A3(KEYINPUT20), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n397_), .A2(new_n398_), .A3(new_n381_), .A4(new_n394_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT101), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT20), .B1(new_n291_), .B2(new_n343_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n343_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n380_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n395_), .A2(new_n400_), .A3(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n404_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT102), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n371_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n404_), .A2(KEYINPUT102), .A3(new_n409_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n409_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n401_), .A2(new_n380_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n336_), .B2(new_n393_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n397_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT97), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n380_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n417_), .B2(new_n380_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n414_), .B(new_n416_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT103), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n420_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(new_n418_), .A3(new_n380_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n426_), .A2(KEYINPUT103), .A3(new_n414_), .A4(new_n416_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n412_), .A2(new_n413_), .A3(new_n423_), .A4(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n409_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n421_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n371_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n370_), .A2(new_n428_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n234_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n245_), .B1(new_n434_), .B2(KEYINPUT100), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n231_), .A2(new_n235_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n435_), .B(new_n436_), .C1(KEYINPUT100), .C2(new_n434_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n438_));
  AND2_X1   g237(.A1(KEYINPUT99), .A2(KEYINPUT33), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n246_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n246_), .A2(new_n438_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n430_), .A2(new_n441_), .A3(new_n421_), .A4(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n414_), .A2(KEYINPUT32), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n404_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n446_), .B(new_n247_), .C1(new_n429_), .C2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n361_), .A2(new_n362_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n367_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n433_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G57gat), .ZN(new_n453_));
  INV_X1    g252(.A(G64gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G57gat), .A2(G64gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT11), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461_));
  INV_X1    g260(.A(G78gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT69), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G78gat), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n463_), .A2(new_n465_), .A3(G71gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(G71gat), .B1(new_n463_), .B2(new_n465_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n455_), .A2(new_n458_), .A3(new_n456_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n461_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n463_), .A2(new_n465_), .ZN(new_n471_));
  INV_X1    g270(.A(G71gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n463_), .A2(new_n465_), .A3(G71gat), .ZN(new_n474_));
  AND4_X1   g273(.A1(new_n461_), .A2(new_n473_), .A3(new_n469_), .A4(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n460_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n468_), .A2(new_n461_), .A3(new_n469_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n469_), .A3(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT70), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n479_), .A3(new_n459_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n482_));
  AND2_X1   g281(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n488_));
  INV_X1    g287(.A(G92gat), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n482_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT8), .ZN(new_n500_));
  XOR2_X1   g299(.A(G85gat), .B(G92gat), .Z(new_n501_));
  OR3_X1    g300(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n493_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT67), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n500_), .B(new_n501_), .C1(new_n505_), .C2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n494_), .A2(new_n502_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n500_), .B1(new_n513_), .B2(new_n501_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n498_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n481_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT64), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n520_), .B(new_n523_), .C1(new_n518_), .C2(new_n517_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n470_), .A2(new_n475_), .A3(new_n460_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n459_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n476_), .A2(KEYINPUT72), .A3(new_n480_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT12), .A4(new_n515_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT73), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT12), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n519_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n519_), .B2(new_n532_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n517_), .B(new_n530_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n524_), .B1(new_n535_), .B2(new_n523_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G120gat), .B(G148gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n524_), .B(new_n543_), .C1(new_n535_), .C2(new_n523_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(KEYINPUT75), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n536_), .A2(new_n546_), .A3(new_n541_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n545_), .A2(KEYINPUT13), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT13), .B1(new_n545_), .B2(new_n547_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G169gat), .B(G197gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G15gat), .B(G22gat), .ZN(new_n554_));
  INV_X1    g353(.A(G1gat), .ZN(new_n555_));
  INV_X1    g354(.A(G8gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G1gat), .B(G8gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G29gat), .B(G36gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n356_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT76), .B(G43gat), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT77), .B(KEYINPUT15), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n563_), .B(new_n564_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n568_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n561_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n570_), .A2(new_n560_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n573_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n570_), .A2(new_n560_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n574_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n553_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n569_), .A2(new_n572_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n574_), .B(new_n578_), .C1(new_n582_), .C2(new_n561_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n580_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n553_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n550_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n452_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n569_), .A2(new_n572_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n515_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT35), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n516_), .A2(new_n567_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n595_), .A2(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n600_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n592_), .A2(new_n608_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n601_), .A2(KEYINPUT78), .A3(new_n607_), .A4(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT78), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(KEYINPUT79), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n601_), .A2(new_n609_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n604_), .A2(new_n605_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n618_), .A3(new_n606_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(KEYINPUT79), .A3(new_n611_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n615_), .A2(new_n619_), .B1(new_n620_), .B2(new_n614_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n560_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n481_), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT81), .B(G127gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(G155gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n628_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n525_), .A3(KEYINPUT17), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n625_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n625_), .B(new_n633_), .C1(KEYINPUT17), .C2(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n590_), .A2(new_n622_), .A3(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n555_), .A3(new_n247_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT104), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n638_), .A2(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(KEYINPUT104), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n619_), .A2(new_n611_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n636_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n452_), .A2(new_n589_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n247_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .A4(new_n649_), .ZN(G1324gat));
  NAND2_X1  g449(.A1(new_n428_), .A2(new_n432_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n637_), .A2(new_n556_), .A3(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n452_), .A2(new_n589_), .A3(new_n651_), .A4(new_n646_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(new_n654_), .A3(G8gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n653_), .B2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT106), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n652_), .B(new_n660_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n658_), .A2(new_n659_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n647_), .B2(new_n367_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT41), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n637_), .A2(new_n302_), .A3(new_n311_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n647_), .B2(new_n450_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  INV_X1    g469(.A(new_n637_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n449_), .A2(new_n345_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT107), .Z(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n671_), .B2(new_n673_), .ZN(G1327gat));
  INV_X1    g473(.A(new_n636_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n644_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT109), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n452_), .A2(new_n589_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT110), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n452_), .A2(new_n680_), .A3(new_n589_), .A4(new_n677_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n247_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n622_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n433_), .B2(new_n451_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n621_), .B(new_n688_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n370_), .A2(new_n428_), .A3(new_n432_), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n311_), .B(new_n449_), .C1(new_n443_), .C2(new_n447_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n687_), .B1(new_n692_), .B2(KEYINPUT43), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n550_), .A2(new_n675_), .A3(new_n588_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n684_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n685_), .B1(new_n452_), .B2(new_n689_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT44), .B(new_n694_), .C1(new_n697_), .C2(new_n687_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n247_), .A2(G29gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n683_), .B1(new_n699_), .B2(new_n700_), .ZN(G1328gat));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n679_), .A2(new_n702_), .A3(new_n651_), .A4(new_n681_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT45), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n696_), .A2(new_n651_), .A3(new_n698_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(new_n706_), .A3(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(G43gat), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n367_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n696_), .A2(new_n698_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT111), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n682_), .A2(new_n311_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n712_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n696_), .A2(new_n718_), .A3(new_n698_), .A4(new_n713_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n715_), .A2(new_n721_), .A3(new_n717_), .A4(new_n719_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1330gat));
  NAND3_X1  g524(.A1(new_n696_), .A2(new_n449_), .A3(new_n698_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n726_), .A2(KEYINPUT113), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(KEYINPUT113), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(G50gat), .A3(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n682_), .A2(new_n356_), .A3(new_n449_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1331gat));
  INV_X1    g530(.A(new_n550_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(new_n587_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n452_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n646_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n735_), .A2(new_n453_), .A3(new_n648_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n621_), .A3(new_n675_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n247_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n736_), .B1(new_n739_), .B2(new_n453_), .ZN(G1332gat));
  INV_X1    g539(.A(new_n651_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G64gat), .B1(new_n735_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT48), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(new_n454_), .A3(new_n651_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n735_), .B2(new_n367_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n738_), .A2(new_n472_), .A3(new_n311_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n735_), .B2(new_n450_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n738_), .A2(new_n462_), .A3(new_n449_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1335gat));
  AND2_X1   g552(.A1(new_n734_), .A2(new_n677_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n247_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n636_), .B(new_n733_), .C1(new_n697_), .C2(new_n687_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n757_));
  INV_X1    g556(.A(new_n687_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n621_), .B(KEYINPUT108), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n433_), .B2(new_n451_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n760_), .B2(new_n685_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n636_), .A4(new_n733_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n648_), .B1(new_n757_), .B2(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n487_), .A2(new_n488_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n755_), .B1(new_n764_), .B2(new_n766_), .ZN(G1336gat));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n489_), .B(new_n741_), .C1(new_n757_), .C2(new_n763_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n734_), .A2(new_n651_), .A3(new_n677_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n489_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n769_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n757_), .A2(new_n763_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(G92gat), .A3(new_n651_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n771_), .B(KEYINPUT115), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(KEYINPUT116), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n778_), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n756_), .B2(new_n367_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n754_), .A2(new_n495_), .A3(new_n311_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n780_), .B(new_n781_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n783_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n754_), .A2(new_n496_), .A3(new_n449_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n761_), .A2(new_n636_), .A3(new_n449_), .A4(new_n733_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(G106gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n788_), .B2(G106gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n787_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1339gat));
  NAND2_X1  g595(.A1(new_n578_), .A2(new_n579_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n574_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n578_), .B1(new_n582_), .B2(new_n561_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n798_), .B(new_n553_), .C1(new_n799_), .C2(new_n574_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(new_n586_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n535_), .A2(new_n523_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT55), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n535_), .A2(new_n523_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n535_), .A2(new_n806_), .A3(new_n523_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n541_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n806_), .B1(new_n535_), .B2(new_n523_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n535_), .A2(new_n523_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT56), .B(new_n541_), .C1(new_n813_), .C2(new_n807_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n544_), .B(new_n801_), .C1(new_n810_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n541_), .B1(new_n813_), .B2(new_n807_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n814_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n822_), .A2(KEYINPUT58), .A3(new_n544_), .A4(new_n801_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n622_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n587_), .A2(new_n544_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT119), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n587_), .A2(new_n544_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n821_), .B2(new_n814_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n545_), .A2(new_n547_), .A3(new_n801_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n644_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT57), .B(new_n644_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n824_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n636_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n587_), .A2(new_n636_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT118), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n621_), .B(new_n839_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n837_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n363_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n651_), .A2(new_n648_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n587_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n588_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n853_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n732_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n848_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n732_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g658(.A(G127gat), .B1(new_n848_), .B2(new_n675_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(G127gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G127gat), .B1(new_n636_), .B2(new_n861_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n860_), .B1(new_n863_), .B2(new_n864_), .ZN(G1342gat));
  AOI21_X1  g664(.A(G134gat), .B1(new_n848_), .B2(new_n645_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n621_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g667(.A(new_n369_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n846_), .A2(new_n869_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT122), .Z(new_n871_));
  AOI21_X1  g670(.A(new_n842_), .B1(new_n836_), .B2(new_n636_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n587_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n550_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n675_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n873_), .B2(new_n645_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n689_), .A2(G162gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n873_), .B2(new_n882_), .ZN(G1347gat));
  NOR3_X1   g682(.A1(new_n872_), .A2(new_n247_), .A3(new_n741_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n845_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n885_), .A2(new_n588_), .A3(new_n288_), .ZN(new_n886_));
  INV_X1    g685(.A(G169gat), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n872_), .A2(new_n247_), .A3(new_n363_), .A4(new_n741_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n587_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT62), .B1(new_n886_), .B2(new_n889_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n889_), .A2(KEYINPUT62), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1348gat));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n550_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n888_), .A2(new_n675_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n385_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n260_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n888_), .A2(KEYINPUT123), .A3(new_n675_), .A4(new_n271_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n885_), .B2(new_n621_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n888_), .A2(new_n645_), .A3(new_n266_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1351gat));
  NAND4_X1  g702(.A1(new_n844_), .A2(new_n648_), .A3(new_n869_), .A4(new_n651_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT124), .B1(new_n884_), .B2(new_n869_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n587_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G197gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n904_), .A2(new_n905_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n872_), .A2(new_n247_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n911_), .A2(KEYINPUT124), .A3(new_n869_), .A4(new_n651_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(G197gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n914_), .A3(new_n587_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n909_), .A2(new_n915_), .ZN(G1352gat));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G204gat), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT126), .Z(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(new_n913_), .B2(new_n550_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n919_), .ZN(new_n921_));
  AOI211_X1 g720(.A(new_n732_), .B(new_n921_), .C1(new_n910_), .C2(new_n912_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n922_), .ZN(G1353gat));
  OR2_X1    g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n913_), .B2(new_n675_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT63), .B(G211gat), .ZN(new_n926_));
  AOI211_X1 g725(.A(new_n636_), .B(new_n926_), .C1(new_n910_), .C2(new_n912_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1354gat));
  NAND2_X1  g727(.A1(new_n913_), .A2(new_n645_), .ZN(new_n929_));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n621_), .A2(new_n930_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT127), .ZN(new_n932_));
  AOI22_X1  g731(.A1(new_n929_), .A2(new_n930_), .B1(new_n913_), .B2(new_n932_), .ZN(G1355gat));
endmodule


