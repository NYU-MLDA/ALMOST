//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XOR2_X1   g001(.A(G8gat), .B(G36gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(G197gat), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G204gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT92), .B1(new_n210_), .B2(G197gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT21), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT92), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n217_), .A3(G197gat), .A4(new_n208_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT21), .B1(new_n213_), .B2(new_n218_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT91), .B(G204gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(G197gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n215_), .B1(G197gat), .B2(G204gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n214_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n219_), .B1(new_n220_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n227_), .A2(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(KEYINPUT24), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT23), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(G183gat), .A3(G190gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT84), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT84), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(new_n238_), .B2(KEYINPUT23), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT22), .B(G169gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT83), .B(G176gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n235_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  OAI22_X1  g049(.A1(new_n237_), .A2(new_n245_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n226_), .A2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n252_), .A2(KEYINPUT20), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n226_), .A2(KEYINPUT93), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT93), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n255_), .B(new_n219_), .C1(new_n220_), .C2(new_n225_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  OAI22_X1  g056(.A1(new_n242_), .A2(new_n244_), .B1(G183gat), .B2(G190gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n235_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT22), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(G169gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n261_), .A2(KEYINPUT82), .B1(G169gat), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n249_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n259_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n239_), .A2(new_n241_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n234_), .A2(KEYINPUT81), .A3(KEYINPUT24), .A4(new_n235_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n236_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n231_), .A2(new_n267_), .A3(new_n268_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n266_), .A2(new_n271_), .A3(KEYINPUT85), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n253_), .B1(new_n257_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n266_), .A2(KEYINPUT85), .A3(new_n271_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT85), .B1(new_n266_), .B2(new_n271_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n254_), .B(new_n256_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n226_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n251_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n280_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n206_), .B1(new_n281_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n252_), .A2(KEYINPUT20), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n282_), .A2(new_n283_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n254_), .A2(new_n256_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n280_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n288_), .B(new_n206_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n202_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT101), .ZN(new_n298_));
  INV_X1    g097(.A(new_n206_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n291_), .A2(new_n292_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n294_), .B1(new_n300_), .B2(new_n253_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n287_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n299_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n295_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT101), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n202_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n298_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n226_), .B(KEYINPUT95), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(new_n251_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n284_), .A2(KEYINPUT20), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n280_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n293_), .A2(new_n294_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n299_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(KEYINPUT27), .A3(new_n295_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G134gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G127gat), .ZN(new_n319_));
  INV_X1    g118(.A(G127gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G134gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n317_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n320_), .A2(G134gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n318_), .A2(G127gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT87), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n319_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n316_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT31), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(G15gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT30), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n332_), .B(new_n336_), .Z(new_n337_));
  XOR2_X1   g136(.A(G71gat), .B(G99gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT86), .B(G43gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n276_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n337_), .B(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT94), .ZN(new_n344_));
  INV_X1    g143(.A(G141gat), .ZN(new_n345_));
  INV_X1    g144(.A(G148gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT3), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT90), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n351_), .A2(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n350_), .B(new_n355_), .C1(new_n352_), .C2(new_n351_), .ZN(new_n356_));
  OR3_X1    g155(.A1(KEYINPUT89), .A2(G155gat), .A3(G162gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(KEYINPUT1), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(G155gat), .A3(G162gat), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n357_), .A2(new_n363_), .A3(new_n365_), .A4(new_n358_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G141gat), .B(G148gat), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n362_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n344_), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n356_), .A2(new_n361_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n371_), .A2(KEYINPUT94), .A3(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n343_), .B1(new_n308_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n369_), .A2(KEYINPUT29), .B1(G228gat), .B2(G233gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n257_), .A2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT28), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n371_), .A2(new_n380_), .A3(new_n372_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n379_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT96), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n379_), .A2(new_n381_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n382_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n392_), .B2(new_n384_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n376_), .B(new_n378_), .C1(new_n388_), .C2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n389_), .B(new_n387_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n387_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n396_), .A3(new_n384_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n378_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n395_), .B(new_n397_), .C1(new_n375_), .C2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n351_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n349_), .A2(new_n347_), .B1(new_n401_), .B2(KEYINPUT90), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n360_), .B1(new_n402_), .B2(new_n355_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n366_), .A2(new_n367_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n331_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n362_), .A2(new_n330_), .A3(new_n325_), .A4(new_n368_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT4), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT98), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT98), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n405_), .A2(new_n406_), .A3(new_n409_), .A4(KEYINPUT4), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT100), .B(KEYINPUT4), .Z(new_n412_));
  NAND3_X1  g211(.A1(new_n369_), .A2(new_n331_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT99), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n405_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n406_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n415_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G85gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT0), .B(G57gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  NAND3_X1  g225(.A1(new_n418_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n426_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n416_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n429_), .B2(new_n421_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n400_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n307_), .A2(new_n315_), .A3(new_n342_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n431_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n400_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n295_), .A2(KEYINPUT27), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(new_n299_), .B2(new_n313_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n427_), .A2(new_n439_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n429_), .A2(new_n421_), .A3(new_n428_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT33), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n415_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n411_), .A2(new_n444_), .A3(new_n413_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n419_), .A2(new_n420_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n426_), .B1(new_n446_), .B2(new_n415_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n303_), .A2(new_n295_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n288_), .B(new_n450_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n426_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n441_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n450_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n443_), .A2(new_n449_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n400_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n307_), .A2(new_n438_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n342_), .B(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n433_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G29gat), .B(G36gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G43gat), .B(G50gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT15), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  INV_X1    g265(.A(G1gat), .ZN(new_n467_));
  INV_X1    g266(.A(G8gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT14), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G8gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n465_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n464_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G229gat), .A2(G233gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n472_), .B(new_n474_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n476_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G113gat), .B(G141gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(KEYINPUT78), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n481_), .A2(KEYINPUT79), .A3(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT80), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n482_), .A2(new_n487_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n490_), .B(new_n491_), .C1(KEYINPUT79), .C2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(KEYINPUT79), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n486_), .A2(new_n489_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT80), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n461_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G232gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT35), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT8), .ZN(new_n505_));
  XOR2_X1   g304(.A(G85gat), .B(G92gat), .Z(new_n506_));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT7), .ZN(new_n508_));
  NOR2_X1   g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n510_), .B1(new_n511_), .B2(new_n509_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT6), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT6), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(G99gat), .A3(G106gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n505_), .B(new_n506_), .C1(new_n512_), .C2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n506_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT67), .B1(new_n514_), .B2(new_n516_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT7), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT66), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n509_), .B1(new_n508_), .B2(new_n523_), .ZN(new_n524_));
  AOI211_X1 g323(.A(G99gat), .B(G106gat), .C1(new_n507_), .C2(KEYINPUT7), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n521_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT67), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n517_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n520_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n519_), .B1(new_n530_), .B2(new_n505_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n506_), .A2(KEYINPUT9), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT65), .B(G85gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT9), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(G92gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n517_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G106gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT10), .B(G99gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT64), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n531_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(KEYINPUT73), .B(new_n504_), .C1(new_n542_), .C2(new_n474_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n502_), .A2(new_n503_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n465_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n504_), .B1(new_n542_), .B2(new_n474_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n543_), .B(new_n544_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n528_), .A2(new_n512_), .A3(new_n521_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT8), .B1(new_n549_), .B2(new_n520_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n540_), .B1(new_n550_), .B2(new_n519_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n551_), .A2(new_n464_), .B1(new_n503_), .B2(new_n502_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n544_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n552_), .B(new_n545_), .C1(KEYINPUT73), .C2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G190gat), .B(G218gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT74), .Z(new_n560_));
  AND3_X1   g359(.A1(new_n548_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n557_), .B(KEYINPUT36), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n548_), .B2(new_n554_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT76), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n548_), .A2(new_n554_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n562_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT76), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n548_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n564_), .A2(KEYINPUT75), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT37), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n565_), .A2(new_n570_), .A3(new_n572_), .A4(KEYINPUT37), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT16), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n472_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT11), .ZN(new_n584_));
  XOR2_X1   g383(.A(G71gat), .B(G78gat), .Z(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(KEYINPUT11), .B2(new_n583_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n582_), .B(new_n588_), .Z(new_n589_));
  OAI21_X1  g388(.A(new_n580_), .B1(new_n589_), .B2(KEYINPUT17), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(KEYINPUT17), .B2(new_n580_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT77), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n591_), .B(new_n593_), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n576_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n588_), .B1(new_n531_), .B2(new_n541_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT12), .B1(new_n597_), .B2(KEYINPUT68), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT68), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n599_), .B(new_n600_), .C1(new_n551_), .C2(new_n588_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n551_), .B2(new_n588_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n598_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT69), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n551_), .A2(new_n588_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n603_), .B1(new_n608_), .B2(new_n597_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT69), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n598_), .A2(new_n601_), .A3(new_n604_), .A4(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G120gat), .B(G148gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n606_), .A2(new_n609_), .A3(new_n611_), .A4(new_n617_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n619_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT71), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT13), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n596_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n499_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  AOI21_X1  g431(.A(G1gat), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n431_), .A3(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n631_), .A2(new_n632_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n561_), .A2(new_n564_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n461_), .A2(new_n594_), .A3(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n497_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT103), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n641_), .B(new_n497_), .C1(new_n623_), .C2(new_n626_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n638_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT104), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(new_n431_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n636_), .B1(new_n645_), .B2(new_n467_), .ZN(G1324gat));
  NAND2_X1  g445(.A1(new_n307_), .A2(new_n315_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n630_), .A2(new_n468_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n643_), .A2(new_n647_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(G8gat), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT39), .B(new_n468_), .C1(new_n643_), .C2(new_n647_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g453(.A1(new_n630_), .A2(new_n334_), .A3(new_n459_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n644_), .A2(new_n459_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n656_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT41), .B1(new_n656_), .B2(G15gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n630_), .A2(new_n660_), .A3(new_n400_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n644_), .B2(new_n400_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n662_), .A2(new_n663_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n594_), .A2(new_n637_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n627_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n499_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n431_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n640_), .A2(new_n642_), .A3(new_n594_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n640_), .A2(KEYINPUT106), .A3(new_n642_), .A4(new_n594_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n574_), .A2(new_n575_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n431_), .B1(new_n394_), .B2(new_n399_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n305_), .B1(new_n304_), .B2(new_n202_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT101), .B(KEYINPUT27), .C1(new_n303_), .C2(new_n295_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n679_), .B(new_n315_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n455_), .A2(new_n456_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n459_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n315_), .B(new_n342_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n432_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n677_), .B(new_n678_), .C1(new_n684_), .C2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT107), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n460_), .A2(new_n690_), .A3(new_n677_), .A4(new_n678_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n678_), .B1(new_n684_), .B2(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT43), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n689_), .A2(new_n691_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n676_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n676_), .A2(new_n694_), .A3(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n431_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n671_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(new_n647_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n669_), .A2(G36gat), .A3(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n647_), .A3(new_n698_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G36gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G36gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI221_X1 g512(.A(new_n706_), .B1(KEYINPUT110), .B2(KEYINPUT46), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1329gat));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n342_), .A2(G43gat), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n699_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  INV_X1    g518(.A(new_n459_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n669_), .B2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n699_), .B2(new_n717_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n718_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n718_), .A2(new_n725_), .A3(new_n721_), .A4(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n670_), .B2(new_n400_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n400_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n700_), .B2(new_n729_), .ZN(G1331gat));
  NAND3_X1  g529(.A1(new_n638_), .A2(new_n498_), .A3(new_n627_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n434_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n460_), .A2(new_n498_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n627_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n596_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT112), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n434_), .A2(G57gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n732_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  OAI21_X1  g538(.A(G64gat), .B1(new_n731_), .B2(new_n703_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n703_), .A2(G64gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n737_), .B2(new_n743_), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n731_), .B2(new_n720_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT49), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n720_), .A2(G71gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n737_), .B2(new_n747_), .ZN(G1334gat));
  OAI21_X1  g547(.A(G78gat), .B1(new_n731_), .B2(new_n456_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT50), .ZN(new_n750_));
  INV_X1    g549(.A(G78gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n736_), .A2(new_n751_), .A3(new_n400_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT114), .ZN(G1335gat));
  OR3_X1    g553(.A1(new_n733_), .A2(new_n734_), .A3(new_n667_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n431_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n734_), .A2(new_n497_), .A3(new_n595_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n694_), .A2(new_n758_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT115), .Z(new_n760_));
  AND2_X1   g559(.A1(new_n431_), .A2(new_n533_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1336gat));
  INV_X1    g561(.A(G92gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n756_), .A2(new_n763_), .A3(new_n647_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n760_), .A2(new_n647_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n763_), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n759_), .B2(new_n720_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n756_), .A2(new_n539_), .A3(new_n342_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n756_), .A2(new_n537_), .A3(new_n400_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n694_), .A2(KEYINPUT116), .A3(new_n400_), .A4(new_n758_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(G106gat), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n759_), .B2(new_n456_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n773_), .A2(new_n774_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n773_), .B2(new_n776_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n771_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n771_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  NAND2_X1  g582(.A1(new_n628_), .A2(new_n498_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n784_), .B(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n497_), .A2(new_n620_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n605_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n598_), .A2(new_n607_), .A3(new_n601_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n603_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n606_), .A2(new_n789_), .A3(new_n611_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n618_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n788_), .B1(new_n795_), .B2(KEYINPUT118), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n618_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n618_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n796_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n619_), .A2(new_n620_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n473_), .A2(new_n475_), .A3(new_n479_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n485_), .B1(new_n478_), .B2(new_n476_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n482_), .A2(new_n485_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n637_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(KEYINPUT57), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n620_), .A2(new_n807_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n798_), .B(new_n617_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n795_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n576_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n814_), .B(KEYINPUT119), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n820_), .A2(KEYINPUT120), .B1(KEYINPUT58), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n678_), .B1(new_n822_), .B2(KEYINPUT58), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n796_), .A2(new_n802_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n637_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n809_), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n810_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n813_), .A2(new_n827_), .A3(new_n830_), .A4(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n787_), .B1(new_n832_), .B2(new_n594_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n685_), .A2(new_n434_), .A3(new_n400_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT122), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n812_), .A2(new_n811_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n831_), .A2(new_n830_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n595_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n838_), .B(new_n834_), .C1(new_n841_), .C2(new_n787_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n836_), .A2(new_n837_), .A3(new_n842_), .A4(new_n497_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT59), .B(new_n834_), .C1(new_n841_), .C2(new_n787_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n498_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n843_), .B1(new_n847_), .B2(new_n837_), .ZN(G1340gat));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n734_), .B2(KEYINPUT60), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n849_), .A2(KEYINPUT60), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n836_), .A2(new_n842_), .A3(new_n850_), .A4(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n734_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n849_), .ZN(G1341gat));
  NAND4_X1  g653(.A1(new_n836_), .A2(new_n320_), .A3(new_n842_), .A4(new_n595_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n594_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n320_), .ZN(G1342gat));
  NAND4_X1  g656(.A1(new_n836_), .A2(new_n318_), .A3(new_n842_), .A4(new_n637_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n576_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n318_), .ZN(G1343gat));
  NAND4_X1  g659(.A1(new_n703_), .A2(new_n431_), .A3(new_n400_), .A4(new_n720_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n833_), .A2(new_n498_), .A3(new_n861_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT123), .B(G141gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1344gat));
  NOR3_X1   g663(.A1(new_n833_), .A2(new_n734_), .A3(new_n861_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n346_), .ZN(G1345gat));
  NOR3_X1   g665(.A1(new_n833_), .A2(new_n594_), .A3(new_n861_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n867_), .B(new_n869_), .ZN(G1346gat));
  NOR2_X1   g669(.A1(new_n833_), .A2(new_n861_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G162gat), .B1(new_n871_), .B2(new_n637_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n678_), .A2(G162gat), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT124), .Z(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n871_), .B2(new_n874_), .ZN(G1347gat));
  NOR3_X1   g674(.A1(new_n703_), .A2(new_n720_), .A3(new_n686_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n497_), .B(new_n876_), .C1(new_n841_), .C2(new_n787_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n877_), .A2(new_n878_), .A3(G169gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n877_), .B2(G169gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n876_), .B1(new_n841_), .B2(new_n787_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n498_), .A2(new_n248_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT125), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n879_), .A2(new_n880_), .B1(new_n881_), .B2(new_n883_), .ZN(G1348gat));
  NOR3_X1   g683(.A1(new_n881_), .A2(new_n233_), .A3(new_n734_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n881_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n627_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n264_), .B2(new_n887_), .ZN(G1349gat));
  INV_X1    g687(.A(G183gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT126), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n886_), .A2(new_n227_), .A3(new_n595_), .A4(new_n890_), .ZN(new_n891_));
  OAI22_X1  g690(.A1(new_n881_), .A2(new_n594_), .B1(KEYINPUT126), .B2(G183gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n881_), .B2(new_n576_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n637_), .A2(new_n228_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n881_), .B2(new_n895_), .ZN(G1351gat));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n703_), .A2(new_n435_), .A3(new_n459_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n497_), .B(new_n898_), .C1(new_n841_), .C2(new_n787_), .ZN(new_n899_));
  INV_X1    g698(.A(G197gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n898_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n832_), .A2(new_n594_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n787_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n905_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n497_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n899_), .A2(new_n900_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n901_), .A2(new_n906_), .A3(new_n907_), .ZN(G1352gat));
  AOI21_X1  g707(.A(G204gat), .B1(new_n905_), .B2(new_n627_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n833_), .A2(new_n734_), .A3(new_n902_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n221_), .B2(new_n910_), .ZN(G1353gat));
  AOI211_X1 g710(.A(KEYINPUT63), .B(G211gat), .C1(new_n905_), .C2(new_n595_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT63), .B(G211gat), .ZN(new_n913_));
  NOR4_X1   g712(.A1(new_n833_), .A2(new_n594_), .A3(new_n902_), .A4(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n912_), .A2(new_n914_), .ZN(G1354gat));
  INV_X1    g714(.A(G218gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n905_), .A2(new_n916_), .A3(new_n637_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n833_), .A2(new_n576_), .A3(new_n902_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n916_), .B2(new_n918_), .ZN(G1355gat));
endmodule


