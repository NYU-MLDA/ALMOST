//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n833_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT93), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  INV_X1    g003(.A(G43gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G50gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(G43gat), .ZN(new_n208_));
  INV_X1    g007(.A(G50gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n207_), .A2(new_n210_), .A3(KEYINPUT15), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216_));
  INV_X1    g015(.A(G1gat), .ZN(new_n217_));
  INV_X1    g016(.A(G8gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G1gat), .B(G8gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n220_), .B(new_n221_), .Z(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n207_), .A3(new_n210_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n211_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n226_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n225_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n223_), .A2(new_n211_), .A3(KEYINPUT75), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(G197gat), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n238_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n227_), .A2(new_n233_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT10), .B(G99gat), .Z(new_n243_));
  INV_X1    g042(.A(G106gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G85gat), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n246_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(KEYINPUT64), .ZN(new_n248_));
  OAI21_X1  g047(.A(G92gat), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n246_), .A2(G92gat), .ZN(new_n254_));
  INV_X1    g053(.A(G92gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(G85gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT9), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n245_), .A2(new_n249_), .A3(new_n253_), .A4(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT8), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G85gat), .B(G92gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT66), .B1(new_n251_), .B2(new_n252_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G99gat), .A2(G106gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT6), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n250_), .ZN(new_n269_));
  OR3_X1    g068(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n263_), .A2(new_n264_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n259_), .B1(new_n262_), .B2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n270_), .A2(new_n264_), .A3(new_n267_), .A4(new_n250_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n260_), .A2(new_n261_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n254_), .A2(new_n256_), .A3(KEYINPUT65), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n259_), .B(new_n273_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n258_), .B1(new_n272_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n281_));
  XOR2_X1   g080(.A(G71gat), .B(G78gat), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n285_), .B(new_n258_), .C1(new_n272_), .C2(new_n277_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G230gat), .A2(G233gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT67), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(KEYINPUT67), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT12), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT68), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n278_), .A2(new_n286_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n278_), .B2(new_n286_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(KEYINPUT68), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n288_), .A2(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n297_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n290_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n293_), .A2(new_n294_), .A3(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G120gat), .B(G148gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G204gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT5), .ZN(new_n306_));
  INV_X1    g105(.A(G176gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT13), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n293_), .A2(new_n302_), .A3(new_n294_), .A4(new_n308_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n242_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT25), .B(G183gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT26), .B(G190gat), .ZN(new_n318_));
  INV_X1    g117(.A(G183gat), .ZN(new_n319_));
  INV_X1    g118(.A(G190gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT23), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(G183gat), .A3(G190gat), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n317_), .A2(new_n318_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT24), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT87), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT24), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(KEYINPUT76), .A2(G169gat), .A3(G176gat), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n326_), .B(new_n328_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n328_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n236_), .A3(new_n307_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n333_), .A2(new_n334_), .A3(new_n336_), .A4(new_n329_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n324_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G169gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n307_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n334_), .B(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n321_), .A2(new_n323_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n340_), .B(new_n342_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT90), .ZN(new_n347_));
  OR2_X1    g146(.A1(G211gat), .A2(G218gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G211gat), .A2(G218gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT84), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT21), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G197gat), .B(G204gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n349_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n351_), .B(new_n353_), .C1(KEYINPUT21), .C2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT90), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n338_), .A2(new_n345_), .A3(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n347_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n330_), .A2(new_n331_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n362_), .A2(new_n342_), .A3(new_n363_), .A4(KEYINPUT24), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n336_), .A2(KEYINPUT24), .A3(new_n329_), .ZN(new_n365_));
  AND3_X1   g164(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT78), .B1(new_n365_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n325_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n364_), .A2(new_n369_), .A3(new_n324_), .A4(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n345_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n357_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n361_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n376_), .B(KEYINPUT86), .Z(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT19), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n346_), .A2(new_n357_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n381_), .B(KEYINPUT20), .C1(new_n372_), .C2(new_n357_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(new_n379_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT18), .B(G64gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G92gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(KEYINPUT32), .A3(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G127gat), .A2(G134gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G113gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G127gat), .A2(G134gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(G127gat), .A2(G134gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(G113gat), .B1(new_n395_), .B2(new_n390_), .ZN(new_n396_));
  AOI21_X1  g195(.A(G120gat), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n396_), .A3(G120gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT81), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n406_), .A3(KEYINPUT2), .ZN(new_n407_));
  AND2_X1   g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT83), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n405_), .B(new_n407_), .C1(new_n410_), .C2(KEYINPUT2), .ZN(new_n411_));
  OR2_X1    g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n403_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n402_), .B2(KEYINPUT1), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n402_), .A2(KEYINPUT1), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n419_), .A2(KEYINPUT82), .A3(G155gat), .A4(G162gat), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n417_), .A2(new_n401_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n409_), .A2(G141gat), .A3(G148gat), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n405_), .A4(new_n412_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n400_), .B1(new_n415_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n403_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT2), .B1(new_n422_), .B2(new_n406_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n405_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n404_), .A2(new_n406_), .A3(KEYINPUT2), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n412_), .B(KEYINPUT3), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n426_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n394_), .A2(new_n396_), .A3(G120gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(new_n397_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n434_), .A3(new_n423_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n425_), .A2(new_n435_), .A3(KEYINPUT4), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n423_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n400_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n425_), .B2(new_n435_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT0), .B(G57gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G85gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(G1gat), .B(G29gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n443_), .A2(new_n445_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n441_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n449_), .B1(new_n452_), .B2(new_n444_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT20), .B1(new_n346_), .B2(new_n357_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n371_), .A2(new_n345_), .B1(new_n356_), .B2(new_n355_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n379_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n346_), .A2(new_n357_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n373_), .A2(new_n460_), .A3(KEYINPUT20), .A4(new_n378_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT88), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n382_), .A2(new_n379_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n388_), .A2(KEYINPUT32), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n459_), .A2(new_n462_), .A3(new_n463_), .A4(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n389_), .A2(new_n454_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n388_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n463_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n461_), .A2(KEYINPUT88), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n453_), .A2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n459_), .A2(new_n462_), .A3(new_n388_), .A4(new_n463_), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT33), .B(new_n449_), .C1(new_n452_), .C2(new_n444_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n470_), .A2(new_n472_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n440_), .A2(new_n442_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n425_), .A2(new_n435_), .A3(new_n442_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n476_), .A2(new_n449_), .A3(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n466_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G22gat), .B(G50gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT28), .ZN(new_n481_));
  OR3_X1    g280(.A1(new_n437_), .A2(KEYINPUT29), .A3(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n481_), .B1(new_n437_), .B2(KEYINPUT29), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT85), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(KEYINPUT85), .A3(new_n483_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n437_), .A2(KEYINPUT29), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n357_), .ZN(new_n488_));
  INV_X1    g287(.A(G228gat), .ZN(new_n489_));
  INV_X1    g288(.A(G233gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n487_), .B(new_n357_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G78gat), .B(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n485_), .B(new_n486_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n484_), .A3(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n479_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT91), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n502_), .A2(new_n454_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n384_), .A2(new_n467_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(KEYINPUT27), .A3(new_n473_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT27), .B1(new_n470_), .B2(new_n473_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n508_), .A2(new_n509_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n505_), .B(new_n507_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n479_), .A2(new_n502_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G227gat), .A2(G233gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT30), .Z(new_n517_));
  XNOR2_X1  g316(.A(new_n434_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G43gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT79), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n518_), .B(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G71gat), .B(G99gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n372_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n523_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n515_), .A2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n507_), .B(new_n502_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n526_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n454_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n316_), .B1(new_n527_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n215_), .A2(new_n278_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n278_), .A2(new_n211_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT69), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n536_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n535_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n540_), .A2(new_n541_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT70), .A4(new_n542_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT71), .B(G134gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G162gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n553_));
  OAI221_X1 g352(.A(new_n535_), .B1(new_n541_), .B2(new_n540_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n548_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n548_), .A2(new_n558_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(KEYINPUT73), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n222_), .B(new_n285_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G183gat), .B(G211gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  OR3_X1    g371(.A1(new_n566_), .A2(new_n567_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(KEYINPUT17), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n566_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n557_), .A2(KEYINPUT73), .A3(KEYINPUT37), .A4(new_n559_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n562_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n203_), .B1(new_n534_), .B2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n532_), .B1(new_n515_), .B2(new_n526_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n562_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n582_));
  NOR4_X1   g381(.A1(new_n581_), .A2(KEYINPUT93), .A3(new_n582_), .A4(new_n316_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n202_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n316_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n479_), .A2(new_n513_), .A3(new_n502_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n513_), .B1(new_n479_), .B2(new_n502_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n529_), .B1(new_n588_), .B2(new_n512_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n585_), .B(new_n579_), .C1(new_n589_), .C2(new_n532_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT93), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n534_), .A2(new_n203_), .A3(new_n579_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(KEYINPUT94), .A3(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n584_), .A2(new_n593_), .A3(new_n217_), .A4(new_n454_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n557_), .A2(new_n559_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n534_), .A2(new_n577_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n530_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n217_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT97), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n603_), .A2(new_n606_), .A3(new_n217_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n596_), .B(new_n597_), .C1(new_n605_), .C2(new_n607_), .ZN(G1324gat));
  OR2_X1    g407(.A1(new_n510_), .A2(new_n511_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n507_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n534_), .A2(new_n577_), .A3(new_n610_), .A4(new_n598_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(G8gat), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT39), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n614_), .A3(G8gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n617_));
  INV_X1    g416(.A(new_n610_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(G8gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n584_), .A2(new_n593_), .A3(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n616_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n617_), .B1(new_n616_), .B2(new_n620_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n584_), .A2(new_n593_), .A3(new_n619_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n611_), .A2(new_n614_), .A3(G8gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n614_), .B1(new_n611_), .B2(G8gat), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT98), .B1(new_n625_), .B2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n616_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT40), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n624_), .A2(new_n631_), .ZN(G1325gat));
  NOR2_X1   g431(.A1(new_n580_), .A2(new_n583_), .ZN(new_n633_));
  INV_X1    g432(.A(G15gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n529_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n601_), .A2(new_n602_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n529_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n637_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT41), .B1(new_n637_), .B2(G15gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(G1326gat));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n502_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n633_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n636_), .A2(new_n642_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(G22gat), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT42), .B(new_n641_), .C1(new_n636_), .C2(new_n642_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(G1327gat));
  NAND2_X1  g447(.A1(new_n585_), .A2(new_n576_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n581_), .A2(new_n649_), .A3(new_n598_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n454_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n562_), .A2(new_n578_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT43), .B1(new_n581_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n655_), .B(new_n652_), .C1(new_n589_), .C2(new_n532_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n649_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(KEYINPUT99), .A3(KEYINPUT44), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n649_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n661_));
  OR2_X1    g460(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n530_), .B1(new_n660_), .B2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n651_), .B1(new_n665_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g465(.A(G36gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n650_), .A2(new_n667_), .A3(new_n610_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT100), .B(KEYINPUT45), .Z(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT101), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n668_), .B(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n618_), .B1(new_n660_), .B2(new_n664_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n667_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(KEYINPUT102), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT102), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n671_), .C1(new_n672_), .C2(new_n667_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1329gat));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AND4_X1   g479(.A1(new_n658_), .A2(new_n657_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n663_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n529_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G43gat), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n650_), .A2(new_n205_), .A3(new_n529_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n680_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n679_), .B(new_n685_), .C1(new_n683_), .C2(G43gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1330gat));
  AOI21_X1  g488(.A(G50gat), .B1(new_n650_), .B2(new_n642_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n209_), .B1(new_n660_), .B2(new_n664_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n642_), .ZN(G1331gat));
  INV_X1    g491(.A(new_n598_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n314_), .A2(new_n315_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n242_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NOR4_X1   g495(.A1(new_n581_), .A2(new_n576_), .A3(new_n693_), .A4(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(G57gat), .A3(new_n454_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT105), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n581_), .A2(new_n582_), .A3(new_n696_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT104), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n530_), .B1(new_n700_), .B2(KEYINPUT104), .ZN(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n699_), .A2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT106), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n697_), .B2(new_n610_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT48), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n700_), .A2(new_n706_), .A3(new_n610_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1333gat));
  INV_X1    g509(.A(G71gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n697_), .B2(new_n529_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT49), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n700_), .A2(new_n711_), .A3(new_n529_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n697_), .B2(new_n642_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT50), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n700_), .A2(new_n716_), .A3(new_n642_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1335gat));
  NAND3_X1  g519(.A1(new_n694_), .A2(new_n576_), .A3(new_n695_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n581_), .A2(new_n598_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n246_), .B1(new_n723_), .B2(new_n530_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n721_), .B(KEYINPUT107), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n246_), .A2(KEYINPUT64), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n454_), .B1(new_n248_), .B2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n724_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT108), .Z(G1336gat));
  AOI21_X1  g530(.A(G92gat), .B1(new_n722_), .B2(new_n610_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n610_), .A2(G92gat), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT109), .Z(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n726_), .B2(new_n734_), .ZN(G1337gat));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(KEYINPUT51), .ZN(new_n737_));
  OAI21_X1  g536(.A(G99gat), .B1(new_n727_), .B2(new_n526_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n722_), .A2(new_n243_), .A3(new_n529_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(KEYINPUT51), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n740_), .B(new_n741_), .Z(G1338gat));
  NAND3_X1  g541(.A1(new_n722_), .A2(new_n244_), .A3(new_n642_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n726_), .A2(new_n642_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(G106gat), .ZN(new_n746_));
  AOI211_X1 g545(.A(KEYINPUT52), .B(new_n244_), .C1(new_n726_), .C2(new_n642_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n752_));
  INV_X1    g551(.A(new_n315_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n242_), .B1(new_n753_), .B2(new_n313_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n579_), .A2(new_n751_), .A3(new_n752_), .A4(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n754_), .A2(new_n562_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(KEYINPUT111), .A3(new_n750_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n242_), .A2(new_n312_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  INV_X1    g559(.A(new_n296_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n287_), .A2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n288_), .A2(new_n299_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n278_), .A2(new_n286_), .A3(new_n296_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n760_), .B1(new_n765_), .B2(new_n291_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n291_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n765_), .A2(new_n760_), .A3(new_n291_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n309_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT56), .B(new_n309_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n759_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n224_), .A2(new_n231_), .A3(new_n226_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n230_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n238_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n241_), .A2(new_n777_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n778_), .A2(KEYINPUT112), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(KEYINPUT112), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n779_), .A2(new_n780_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n598_), .B1(new_n774_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT113), .B(new_n598_), .C1(new_n774_), .C2(new_n781_), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n786_));
  NAND3_X1  g585(.A1(new_n784_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT55), .B1(new_n301_), .B2(new_n290_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n302_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n769_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n771_), .B(new_n308_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n791_), .A2(KEYINPUT115), .B1(new_n779_), .B2(new_n780_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n772_), .A2(new_n793_), .A3(new_n773_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n794_), .A3(new_n312_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n792_), .A2(new_n794_), .A3(KEYINPUT58), .A4(new_n312_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n652_), .A3(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT57), .B(new_n598_), .C1(new_n774_), .C2(new_n781_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n787_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n758_), .B1(new_n801_), .B2(new_n576_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n642_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n610_), .A2(new_n530_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(new_n526_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n242_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n803_), .A2(KEYINPUT59), .A3(new_n806_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n695_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n809_), .B1(new_n813_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  INV_X1    g614(.A(new_n694_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(KEYINPUT60), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n808_), .B(new_n817_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n815_), .ZN(G1341gat));
  AOI21_X1  g619(.A(G127gat), .B1(new_n808_), .B2(new_n577_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n576_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g622(.A(G134gat), .B1(new_n808_), .B2(new_n693_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n811_), .A2(new_n812_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT116), .B(G134gat), .Z(new_n826_));
  NOR2_X1   g625(.A1(new_n653_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n825_), .B2(new_n827_), .ZN(G1343gat));
  NOR4_X1   g627(.A1(new_n802_), .A2(new_n529_), .A3(new_n502_), .A4(new_n805_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n242_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT117), .B(G141gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1344gat));
  NAND2_X1  g631(.A1(new_n829_), .A2(new_n694_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n577_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT61), .B(G155gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1346gat));
  AOI21_X1  g636(.A(G162gat), .B1(new_n829_), .B2(new_n693_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n652_), .A2(G162gat), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT118), .Z(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n829_), .B2(new_n840_), .ZN(G1347gat));
  NAND2_X1  g640(.A1(new_n801_), .A2(new_n576_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n758_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n502_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n610_), .A2(new_n530_), .A3(new_n529_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT119), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n845_), .A2(new_n695_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n339_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n848_), .B2(new_n236_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n851_), .A3(new_n853_), .ZN(G1348gat));
  NOR2_X1   g653(.A1(new_n845_), .A2(new_n847_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G176gat), .B1(new_n855_), .B2(new_n694_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n803_), .A2(KEYINPUT120), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n802_), .B2(new_n642_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n307_), .B(new_n847_), .C1(new_n857_), .C2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n856_), .B1(new_n860_), .B2(new_n694_), .ZN(G1349gat));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n859_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n847_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n577_), .A3(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n576_), .A2(new_n317_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n864_), .A2(new_n319_), .B1(new_n855_), .B2(new_n865_), .ZN(G1350gat));
  NAND4_X1  g665(.A1(new_n803_), .A2(new_n318_), .A3(new_n693_), .A4(new_n863_), .ZN(new_n867_));
  NOR4_X1   g666(.A1(new_n802_), .A2(new_n642_), .A3(new_n653_), .A4(new_n847_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n320_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT121), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n867_), .B(new_n871_), .C1(new_n320_), .C2(new_n868_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(G1351gat));
  XNOR2_X1  g672(.A(KEYINPUT124), .B(G197gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n642_), .A2(new_n530_), .A3(new_n526_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n610_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n876_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n844_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n879_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(KEYINPUT123), .A3(new_n878_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n874_), .B1(new_n886_), .B2(new_n242_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT123), .B1(new_n884_), .B2(new_n878_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n802_), .A2(new_n881_), .A3(new_n877_), .A4(new_n883_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n242_), .B(new_n874_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n891_), .ZN(G1352gat));
  NOR2_X1   g691(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n893_));
  AND2_X1   g692(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n894_));
  OAI221_X1 g693(.A(new_n694_), .B1(new_n893_), .B2(new_n894_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n816_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n893_), .ZN(G1353gat));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT126), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT127), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n900_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n576_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n886_), .A2(new_n902_), .A3(new_n903_), .A4(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n903_), .B(new_n904_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n901_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1354gat));
  AOI21_X1  g707(.A(G218gat), .B1(new_n886_), .B2(new_n693_), .ZN(new_n909_));
  OAI211_X1 g708(.A(G218gat), .B(new_n652_), .C1(new_n888_), .C2(new_n889_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1355gat));
endmodule


