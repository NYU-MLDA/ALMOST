//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT88), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT88), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n210_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT79), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(G169gat), .B2(G176gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n228_), .A3(KEYINPUT89), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT89), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n213_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n217_), .A2(KEYINPUT88), .A3(new_n218_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n209_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AND4_X1   g032(.A1(KEYINPUT24), .A2(new_n223_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n230_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT23), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n236_), .A2(KEYINPUT23), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n239_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n226_), .A2(KEYINPUT24), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n229_), .A2(new_n235_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n244_), .A2(KEYINPUT21), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(KEYINPUT21), .ZN(new_n246_));
  XOR2_X1   g045(.A(G197gat), .B(G204gat), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n246_), .A2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n237_), .B1(G183gat), .B2(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n227_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT22), .B(G169gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(new_n222_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n243_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n240_), .A2(new_n238_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n238_), .B2(new_n237_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n255_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n210_), .B1(new_n212_), .B2(new_n211_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n242_), .A2(new_n237_), .A3(new_n228_), .A4(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n250_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AND4_X1   g067(.A1(KEYINPUT20), .A2(new_n257_), .A3(new_n265_), .A4(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n243_), .A2(new_n256_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n250_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT90), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n251_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n273_), .A2(KEYINPUT20), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(new_n275_), .A3(new_n250_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  AOI211_X1 g076(.A(new_n206_), .B(new_n269_), .C1(new_n277_), .C2(new_n267_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n251_), .B1(new_n243_), .B2(new_n256_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT90), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT95), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n268_), .A4(new_n274_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n272_), .A2(new_n268_), .A3(new_n274_), .A4(new_n276_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT95), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n257_), .A2(new_n265_), .A3(KEYINPUT20), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n267_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n278_), .B1(new_n287_), .B2(new_n206_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT27), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290_));
  INV_X1    g089(.A(new_n206_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n277_), .A2(new_n267_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n269_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n290_), .B1(new_n294_), .B2(new_n278_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298_));
  INV_X1    g097(.A(G141gat), .ZN(new_n299_));
  INV_X1    g098(.A(G148gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n304_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT1), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n312_), .A3(new_n309_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n314_), .A2(new_n302_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n299_), .A2(new_n300_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n250_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(G228gat), .A3(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n311_), .A2(KEYINPUT82), .A3(new_n317_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n250_), .B1(new_n326_), .B2(KEYINPUT83), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G228gat), .A2(G233gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n311_), .A2(KEYINPUT82), .A3(new_n317_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT82), .B1(new_n311_), .B2(new_n317_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT29), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n328_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n322_), .B1(new_n327_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT84), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT85), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n322_), .B(new_n337_), .C1(new_n327_), .C2(new_n333_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(KEYINPUT86), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT86), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n334_), .A2(new_n342_), .A3(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n324_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G22gat), .B(G50gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT28), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n345_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n334_), .A2(new_n336_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n349_), .B1(new_n351_), .B2(new_n340_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n297_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n348_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n355_), .A2(KEYINPUT87), .A3(new_n352_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n296_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n264_), .B(KEYINPUT30), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(G127gat), .A2(G134gat), .ZN(new_n362_));
  INV_X1    g161(.A(G113gat), .ZN(new_n363_));
  INV_X1    g162(.A(G120gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G127gat), .A2(G134gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G113gat), .A2(G120gat), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n367_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n369_), .A3(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT31), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n361_), .B(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G15gat), .B(G43gat), .Z(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n377_), .B(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n375_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT92), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n385_), .B(new_n375_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n373_), .A2(new_n368_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n319_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n384_), .A2(KEYINPUT4), .A3(new_n386_), .A4(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT93), .ZN(new_n390_));
  INV_X1    g189(.A(new_n383_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n383_), .A2(KEYINPUT92), .B1(new_n387_), .B2(new_n319_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n397_), .A2(new_n390_), .A3(KEYINPUT4), .A4(new_n386_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n386_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n395_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G57gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G85gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(G1gat), .B(G29gat), .Z(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n399_), .A2(new_n406_), .A3(new_n401_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n382_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n358_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n294_), .A2(new_n278_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n408_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n394_), .A2(new_n398_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n395_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n418_), .B(new_n406_), .C1(new_n395_), .C2(new_n400_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n402_), .B(new_n407_), .C1(KEYINPUT94), .C2(KEYINPUT33), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n414_), .A2(new_n416_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n291_), .A2(KEYINPUT32), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n287_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n292_), .A2(new_n293_), .A3(new_n422_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n410_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n357_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n357_), .A3(KEYINPUT96), .ZN(new_n431_));
  INV_X1    g230(.A(new_n356_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT87), .B1(new_n355_), .B2(new_n352_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n296_), .A2(new_n411_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n430_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n382_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n413_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n439_));
  XOR2_X1   g238(.A(G120gat), .B(G148gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT72), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G176gat), .B(G204gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G85gat), .B(G92gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT9), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT10), .B(G99gat), .Z(new_n450_));
  INV_X1    g249(.A(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(G85gat), .A3(G92gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT6), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n449_), .A2(new_n452_), .A3(new_n453_), .A4(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n447_), .B(KEYINPUT64), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT7), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n455_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n457_), .A2(new_n458_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n462_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT65), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(KEYINPUT65), .A3(new_n462_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n455_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n458_), .B1(new_n469_), .B2(new_n457_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT67), .B1(new_n464_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n464_), .A2(new_n470_), .A3(KEYINPUT67), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n456_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT66), .B(G71gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G78gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(G57gat), .B(G64gat), .Z(new_n477_));
  INV_X1    g276(.A(KEYINPUT11), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n478_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G78gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n475_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n479_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT68), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n474_), .A2(new_n488_), .A3(KEYINPUT12), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n486_), .B(new_n456_), .C1(new_n470_), .C2(new_n464_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G230gat), .A2(G233gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(KEYINPUT69), .A3(new_n491_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n486_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n464_), .A2(new_n470_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n456_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n489_), .A2(new_n496_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT70), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT70), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n489_), .A2(new_n496_), .A3(new_n505_), .A4(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n491_), .B1(new_n500_), .B2(new_n490_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n446_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  AOI211_X1 g309(.A(new_n508_), .B(new_n445_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n439_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n500_), .A2(new_n501_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n498_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n471_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n487_), .B1(new_n516_), .B2(new_n456_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n513_), .B1(new_n517_), .B2(KEYINPUT12), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n505_), .B1(new_n518_), .B2(new_n496_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n506_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n509_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n445_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n507_), .A2(new_n509_), .A3(new_n446_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(KEYINPUT73), .A3(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n512_), .A2(new_n524_), .A3(KEYINPUT13), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT13), .B1(new_n512_), .B2(new_n524_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT78), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G29gat), .B(G36gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(G43gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G50gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT76), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533_));
  INV_X1    g332(.A(G1gat), .ZN(new_n534_));
  INV_X1    g333(.A(G8gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G1gat), .B(G8gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n531_), .A2(KEYINPUT76), .ZN(new_n541_));
  INV_X1    g340(.A(new_n539_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n531_), .A2(KEYINPUT76), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n531_), .A2(KEYINPUT15), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n531_), .A2(KEYINPUT15), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n539_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT77), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n553_), .B(new_n539_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n552_), .A2(new_n554_), .A3(new_n546_), .A4(new_n544_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n221_), .ZN(new_n557_));
  INV_X1    g356(.A(G197gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n548_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n548_), .B2(new_n555_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n528_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n548_), .A2(new_n555_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n559_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n548_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(KEYINPUT78), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n527_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT16), .B(G183gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G211gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(KEYINPUT68), .A3(KEYINPUT17), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(KEYINPUT17), .B2(new_n573_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n486_), .B(new_n542_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  MUX2_X1   g377(.A(new_n575_), .B(new_n574_), .S(new_n578_), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n438_), .A2(new_n569_), .A3(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n474_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n531_), .B(new_n456_), .C1(new_n470_), .C2(new_n464_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n582_), .B(new_n583_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n585_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n586_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G134gat), .ZN(new_n597_));
  INV_X1    g396(.A(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n594_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(KEYINPUT36), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(KEYINPUT37), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n601_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n600_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n581_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n534_), .A3(new_n410_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT38), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n581_), .A2(new_n608_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT97), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT97), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n411_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n534_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n618_), .A2(KEYINPUT98), .A3(new_n534_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n614_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT99), .ZN(G1324gat));
  NOR3_X1   g423(.A1(new_n611_), .A2(G8gat), .A3(new_n296_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n626_), .B1(new_n615_), .B2(new_n296_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n289_), .A2(new_n295_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n581_), .A2(KEYINPUT100), .A3(new_n608_), .A4(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(G8gat), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT39), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n627_), .A2(new_n632_), .A3(G8gat), .A4(new_n629_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n625_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AOI211_X1 g435(.A(KEYINPUT101), .B(new_n625_), .C1(new_n631_), .C2(new_n633_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  OR3_X1    g440(.A1(new_n611_), .A2(G15gat), .A3(new_n437_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n616_), .A2(new_n617_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n382_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(new_n644_), .B2(G15gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(G1326gat));
  INV_X1    g446(.A(G22gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n612_), .A2(new_n648_), .A3(new_n434_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n643_), .A2(new_n434_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(G22gat), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT42), .B(new_n648_), .C1(new_n643_), .C2(new_n434_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(G1327gat));
  NOR2_X1   g453(.A1(new_n569_), .A2(new_n579_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n427_), .A2(KEYINPUT96), .A3(new_n357_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT96), .B1(new_n427_), .B2(new_n357_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n411_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n628_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n661_), .A2(new_n382_), .B1(new_n358_), .B2(new_n412_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n607_), .A2(new_n600_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n603_), .B1(new_n663_), .B2(KEYINPUT37), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n656_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n438_), .A2(KEYINPUT43), .A3(new_n610_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n655_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n655_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n410_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n672_), .A2(KEYINPUT102), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(KEYINPUT102), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(G29gat), .A3(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n438_), .A2(new_n608_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n655_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n411_), .A2(G29gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(G1328gat));
  NAND3_X1  g478(.A1(new_n669_), .A2(new_n628_), .A3(new_n670_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT103), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n669_), .A2(new_n682_), .A3(new_n628_), .A4(new_n670_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(G36gat), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT104), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n681_), .A2(new_n686_), .A3(G36gat), .A4(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n677_), .A2(G36gat), .A3(new_n296_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT45), .Z(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(KEYINPUT46), .A3(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1329gat));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n677_), .A2(G43gat), .A3(new_n437_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n671_), .A2(new_n382_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(G43gat), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n699_), .A2(new_n700_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n696_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n703_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(KEYINPUT47), .A3(new_n701_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1330gat));
  NAND2_X1  g506(.A1(new_n671_), .A2(new_n434_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT106), .ZN(new_n709_));
  INV_X1    g508(.A(G50gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n434_), .A2(new_n710_), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n709_), .A2(new_n710_), .B1(new_n677_), .B2(new_n711_), .ZN(G1331gat));
  INV_X1    g511(.A(new_n527_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n568_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n715_), .A2(new_n438_), .A3(new_n580_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n610_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n410_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n608_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n411_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(G57gat), .B2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n720_), .B2(new_n296_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n296_), .A2(G64gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n717_), .B2(new_n725_), .ZN(G1333gat));
  OR3_X1    g525(.A1(new_n717_), .A2(G71gat), .A3(new_n437_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n716_), .A2(new_n608_), .A3(new_n382_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G71gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G71gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT107), .Z(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n720_), .B2(new_n357_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n718_), .A2(new_n483_), .A3(new_n434_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n715_), .A2(new_n579_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(new_n676_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n410_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n665_), .A2(new_n666_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n741_), .A2(new_n579_), .A3(new_n715_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(new_n410_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n740_), .B1(new_n743_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g543(.A(G92gat), .B1(new_n739_), .B2(new_n628_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n628_), .A2(G92gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n742_), .B2(new_n746_), .ZN(G1337gat));
  NAND3_X1  g546(.A1(new_n739_), .A2(new_n450_), .A3(new_n382_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n742_), .A2(new_n382_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n749_), .A2(KEYINPUT108), .A3(G99gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT108), .B1(new_n749_), .B2(G99gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n752_), .B(new_n753_), .Z(G1338gat));
  NAND3_X1  g553(.A1(new_n739_), .A2(new_n451_), .A3(new_n434_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n742_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G106gat), .B1(new_n756_), .B2(new_n357_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(KEYINPUT52), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(KEYINPUT52), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g560(.A(new_n560_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT114), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n552_), .A2(new_n544_), .A3(new_n554_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n546_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n566_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n518_), .A2(KEYINPUT55), .A3(new_n496_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n518_), .A2(new_n490_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(G230gat), .A3(G233gat), .ZN(new_n770_));
  INV_X1    g569(.A(new_n507_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n768_), .B(new_n770_), .C1(new_n771_), .C2(KEYINPUT55), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n445_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT56), .B1(new_n772_), .B2(new_n445_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n523_), .B(new_n767_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n775_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n511_), .B1(new_n780_), .B2(new_n773_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n778_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n767_), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n783_), .A3(new_n664_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n568_), .A2(new_n523_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n780_), .B2(new_n773_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n766_), .B1(new_n512_), .B2(new_n524_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n608_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT57), .B(new_n608_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n784_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(new_n580_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n563_), .A2(new_n567_), .A3(new_n579_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT110), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n527_), .A2(KEYINPUT111), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT13), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n510_), .A2(new_n511_), .A3(new_n439_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT73), .B1(new_n522_), .B2(new_n523_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n512_), .A2(new_n524_), .A3(KEYINPUT13), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n664_), .B1(new_n797_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n794_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT111), .B1(new_n527_), .B2(new_n796_), .ZN(new_n809_));
  AND4_X1   g608(.A1(KEYINPUT111), .A2(new_n796_), .A3(new_n801_), .A4(new_n802_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n610_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT113), .A3(KEYINPUT54), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n807_), .B(new_n610_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT112), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n806_), .A2(new_n816_), .A3(new_n807_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n793_), .B1(new_n813_), .B2(new_n818_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n358_), .A2(new_n411_), .A3(new_n437_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n792_), .A2(new_n580_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT116), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n792_), .A2(new_n826_), .A3(new_n580_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n812_), .A2(new_n808_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n823_), .B(new_n820_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n822_), .A2(new_n830_), .A3(new_n568_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G113gat), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n819_), .A2(new_n821_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n363_), .A3(new_n568_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n837_), .A3(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1340gat));
  NAND3_X1  g638(.A1(new_n822_), .A2(new_n830_), .A3(new_n713_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n364_), .B1(new_n527_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n833_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n364_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n841_), .A2(KEYINPUT118), .A3(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1341gat));
  AOI21_X1  g647(.A(G127gat), .B1(new_n833_), .B2(new_n579_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n822_), .A2(new_n830_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n850_), .A2(new_n579_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n851_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g651(.A(G134gat), .B1(new_n833_), .B2(new_n663_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT119), .B(G134gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n610_), .A2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT120), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n850_), .B2(new_n856_), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n819_), .A2(new_n382_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n628_), .A2(new_n357_), .A3(new_n411_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n714_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n299_), .ZN(G1344gat));
  INV_X1    g661(.A(new_n860_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n713_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT121), .B(G148gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1345gat));
  NOR2_X1   g665(.A1(new_n860_), .A2(new_n580_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT61), .B(G155gat), .Z(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT122), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n867_), .B(new_n869_), .ZN(G1346gat));
  NOR3_X1   g669(.A1(new_n860_), .A2(new_n598_), .A3(new_n610_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n863_), .A2(new_n663_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n598_), .B2(new_n872_), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n412_), .A2(new_n296_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n357_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n827_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n826_), .B1(new_n792_), .B2(new_n580_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n813_), .A2(new_n818_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n221_), .B1(new_n880_), .B2(new_n568_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT124), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(KEYINPUT123), .A3(new_n882_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885_));
  INV_X1    g684(.A(new_n875_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n568_), .B(new_n886_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G169gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n885_), .B1(new_n888_), .B2(KEYINPUT62), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n890_), .A3(KEYINPUT62), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n883_), .A2(new_n884_), .A3(new_n889_), .A4(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n880_), .A2(new_n568_), .A3(new_n254_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1348gat));
  AOI21_X1  g693(.A(G176gat), .B1(new_n880_), .B2(new_n713_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n819_), .A2(new_n434_), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n527_), .A2(new_n222_), .A3(new_n296_), .A4(new_n412_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1349gat));
  INV_X1    g697(.A(new_n880_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n899_), .A2(new_n580_), .A3(new_n210_), .ZN(new_n900_));
  INV_X1    g699(.A(G183gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n896_), .A2(new_n579_), .A3(new_n874_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n899_), .B2(new_n610_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n880_), .B1(new_n219_), .B2(new_n214_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n608_), .ZN(G1351gat));
  NOR2_X1   g705(.A1(new_n296_), .A2(new_n659_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n437_), .B(new_n907_), .C1(new_n829_), .C2(new_n793_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n714_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n558_), .ZN(G1352gat));
  INV_X1    g709(.A(new_n908_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n713_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g712(.A1(new_n908_), .A2(new_n580_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT63), .ZN(new_n916_));
  INV_X1    g715(.A(G211gat), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n914_), .A2(new_n915_), .A3(new_n919_), .A4(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n908_), .B2(new_n580_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT125), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n908_), .A2(new_n580_), .A3(new_n918_), .A4(new_n920_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n922_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT126), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n922_), .B(new_n928_), .C1(new_n924_), .C2(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1354gat));
  AOI21_X1  g729(.A(KEYINPUT127), .B1(new_n911_), .B2(new_n663_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n908_), .A2(new_n932_), .A3(new_n608_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(G218gat), .A3(new_n933_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n664_), .A2(G218gat), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n911_), .B2(new_n935_), .ZN(G1355gat));
endmodule


