//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_;
  XNOR2_X1  g000(.A(G57gat), .B(G85gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G1gat), .B(G29gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT90), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT90), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT92), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n210_), .A2(new_n214_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT3), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n217_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT92), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n211_), .A2(new_n213_), .A3(new_n223_), .A4(new_n214_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n216_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n211_), .A2(new_n213_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n227_), .B(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n231_), .B2(new_n226_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n220_), .B(KEYINPUT91), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n225_), .A2(new_n228_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n236_));
  INV_X1    g035(.A(G113gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(G120gat), .ZN(new_n238_));
  INV_X1    g037(.A(G120gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(G113gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G127gat), .A2(G134gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(G127gat), .A2(G134gat), .ZN(new_n242_));
  OAI22_X1  g041(.A1(new_n238_), .A2(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(G127gat), .A2(G134gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(G113gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(G120gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G127gat), .A2(G134gat), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n243_), .A2(KEYINPUT88), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT88), .B1(new_n243_), .B2(new_n248_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n235_), .A2(new_n236_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n225_), .A2(new_n228_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n232_), .A2(new_n233_), .ZN(new_n254_));
  AND4_X1   g053(.A1(new_n248_), .A2(new_n253_), .A3(new_n243_), .A4(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT102), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT102), .B1(new_n235_), .B2(new_n251_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(new_n255_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n209_), .B(new_n252_), .C1(new_n259_), .C2(new_n236_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n257_), .B(new_n208_), .C1(new_n258_), .C2(new_n255_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n207_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n261_), .A3(new_n207_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G228gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n266_), .A2(G228gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(G233gat), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT29), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G211gat), .A2(G218gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G211gat), .A2(G218gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT95), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(G211gat), .A2(G218gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT95), .B1(new_n279_), .B2(new_n274_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT94), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(KEYINPUT21), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(KEYINPUT21), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n277_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n279_), .A2(KEYINPUT95), .A3(new_n274_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT21), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n285_), .A2(new_n288_), .A3(KEYINPUT94), .A4(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n284_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n271_), .B1(new_n273_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n284_), .A2(new_n291_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(new_n270_), .C1(new_n234_), .C2(new_n272_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G78gat), .B(G106gat), .Z(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT28), .B(G22gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n253_), .A2(new_n272_), .A3(new_n254_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(G50gat), .ZN(new_n301_));
  INV_X1    g100(.A(G50gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n234_), .B2(new_n272_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n299_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(G50gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n234_), .A2(new_n272_), .A3(new_n302_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n298_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n297_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n296_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT97), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n301_), .A2(new_n303_), .A3(new_n299_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n298_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT97), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n293_), .A2(new_n295_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n296_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n313_), .A2(new_n314_), .A3(new_n317_), .A4(new_n297_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n310_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G183gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT85), .B1(new_n320_), .B2(KEYINPUT25), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT26), .B(G190gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT25), .B(G183gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n322_), .C1(new_n323_), .C2(KEYINPUT85), .ZN(new_n324_));
  INV_X1    g123(.A(G190gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT23), .B1(new_n320_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(G183gat), .A3(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G169gat), .ZN(new_n330_));
  INV_X1    g129(.A(G176gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT24), .A3(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n332_), .A2(KEYINPUT24), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n324_), .A2(new_n329_), .A3(new_n334_), .A4(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n326_), .A2(new_n328_), .A3(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n327_), .A2(KEYINPUT86), .A3(G183gat), .A4(G190gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n333_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT22), .B(G169gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(new_n331_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n336_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT89), .B1(new_n249_), .B2(new_n250_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT87), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n349_));
  AND4_X1   g148(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n245_), .A2(new_n246_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n243_), .A2(KEYINPUT88), .A3(new_n248_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n347_), .A2(new_n348_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n348_), .B1(new_n347_), .B2(new_n355_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n346_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT89), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT87), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n346_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n347_), .A2(new_n355_), .A3(new_n348_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G15gat), .B(G43gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT31), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n358_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n358_), .B2(new_n364_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT30), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n368_), .A2(new_n369_), .A3(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n356_), .A2(new_n357_), .A3(new_n346_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n362_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n366_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n358_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n373_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n317_), .A2(KEYINPUT96), .A3(new_n297_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n313_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n297_), .A2(KEYINPUT96), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n319_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n374_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n378_), .A2(new_n373_), .A3(new_n379_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n385_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n310_), .A2(new_n318_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n265_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT27), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT20), .B1(new_n294_), .B2(new_n346_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT98), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n329_), .A2(new_n339_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT100), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT100), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n329_), .A2(new_n402_), .A3(new_n339_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n344_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n323_), .A2(new_n322_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n334_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT99), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n335_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n340_), .B(new_n338_), .C1(new_n406_), .C2(KEYINPUT99), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n404_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n294_), .ZN(new_n411_));
  OAI211_X1 g210(.A(KEYINPUT98), .B(KEYINPUT20), .C1(new_n294_), .C2(new_n346_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n397_), .A2(new_n399_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n294_), .A2(new_n346_), .ZN(new_n414_));
  OAI211_X1 g213(.A(KEYINPUT20), .B(new_n414_), .C1(new_n410_), .C2(new_n294_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n399_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n394_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT105), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n415_), .A2(new_n399_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n397_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(new_n399_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n423_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n425_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n426_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n418_), .A2(new_n424_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n413_), .A2(new_n417_), .A3(new_n423_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT27), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n431_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(KEYINPUT104), .A2(KEYINPUT33), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n264_), .A2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n433_), .A2(new_n434_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT104), .B(KEYINPUT33), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n260_), .A2(new_n261_), .A3(new_n207_), .A4(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n259_), .A2(new_n208_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n252_), .B1(new_n259_), .B2(new_n236_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n442_), .B(new_n206_), .C1(new_n443_), .C2(new_n209_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .A4(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT32), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n418_), .B1(new_n446_), .B2(new_n423_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n429_), .A2(KEYINPUT32), .A3(new_n424_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n260_), .A2(new_n261_), .A3(new_n207_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n447_), .B(new_n448_), .C1(new_n449_), .C2(new_n262_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n445_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n319_), .A2(new_n385_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(new_n381_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n393_), .A2(new_n436_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT77), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(G50gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(G50gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT74), .B(G43gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n457_), .A2(new_n460_), .A3(new_n458_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n462_), .A2(KEYINPUT15), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT15), .B1(new_n462_), .B2(new_n463_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT10), .B(G99gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(G99gat), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n471_), .A2(KEYINPUT10), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(KEYINPUT10), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT65), .B(new_n470_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G85gat), .B(G92gat), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT9), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n478_));
  AND3_X1   g277(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(KEYINPUT66), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(G85gat), .ZN(new_n488_));
  INV_X1    g287(.A(G92gat), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT9), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n475_), .A2(new_n477_), .A3(new_n487_), .A4(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n492_));
  NOR2_X1   g291(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n493_));
  OAI22_X1  g292(.A1(new_n492_), .A2(new_n493_), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n479_), .A2(new_n480_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n471_), .A3(new_n470_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n476_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT8), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT8), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n476_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n481_), .A2(new_n486_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n494_), .A2(new_n497_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT70), .B1(new_n500_), .B2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n494_), .A2(new_n497_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n502_), .B1(new_n508_), .B2(new_n487_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n501_), .B1(new_n498_), .B2(new_n476_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n491_), .B1(new_n507_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n466_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT76), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n491_), .B1(new_n510_), .B2(new_n509_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n457_), .A2(new_n460_), .A3(new_n458_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n460_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n514_), .A2(new_n515_), .A3(new_n521_), .A4(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n464_), .A2(new_n465_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n491_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n500_), .A2(new_n506_), .A3(KEYINPUT70), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n511_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n521_), .B(new_n527_), .C1(new_n529_), .C2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT76), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n529_), .A2(new_n533_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n521_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n525_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n528_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540_));
  INV_X1    g339(.A(G162gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT75), .B(G134gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n544_), .B(KEYINPUT36), .Z(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(KEYINPUT36), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n528_), .A2(new_n535_), .A3(new_n538_), .A4(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n455_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n548_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(KEYINPUT77), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT37), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n546_), .A2(KEYINPUT78), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT78), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n553_), .B(new_n548_), .C1(new_n554_), .C2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(G57gat), .A2(G64gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(G57gat), .A2(G64gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT11), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT68), .ZN(new_n565_));
  INV_X1    g364(.A(G71gat), .ZN(new_n566_));
  INV_X1    g365(.A(G78gat), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n561_), .A2(new_n562_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n567_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G57gat), .B(G64gat), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n569_), .B(new_n571_), .C1(new_n572_), .C2(KEYINPUT11), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(KEYINPUT68), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n564_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(KEYINPUT68), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n561_), .A2(new_n562_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n577_), .A2(new_n565_), .A3(new_n569_), .A4(new_n571_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n578_), .A3(new_n563_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G15gat), .B(G22gat), .ZN(new_n581_));
  INV_X1    g380(.A(G1gat), .ZN(new_n582_));
  INV_X1    g381(.A(G8gat), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT14), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G1gat), .B(G8gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n585_), .B(new_n586_), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n580_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT79), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(KEYINPUT79), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n593_));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT17), .A4(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n597_), .B(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n590_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n454_), .A2(new_n558_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT13), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(G204gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT5), .B(G176gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT12), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n531_), .A2(new_n532_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n611_), .B2(new_n491_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n579_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n563_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT71), .B1(new_n612_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT71), .ZN(new_n617_));
  NOR4_X1   g416(.A1(new_n533_), .A2(new_n617_), .A3(new_n610_), .A4(new_n580_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n610_), .B1(new_n517_), .B2(new_n580_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n517_), .A2(new_n580_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n616_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT64), .Z(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(KEYINPUT72), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n513_), .A2(KEYINPUT12), .A3(new_n615_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n617_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n615_), .A2(new_n516_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n615_), .A2(new_n516_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n610_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n612_), .A2(KEYINPUT71), .A3(new_n615_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n628_), .A2(new_n625_), .A3(new_n631_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT72), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n626_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n620_), .A2(new_n630_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT69), .B1(new_n637_), .B2(new_n624_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT69), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n639_), .B(new_n625_), .C1(new_n620_), .C2(new_n630_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n609_), .B1(new_n636_), .B2(new_n642_), .ZN(new_n643_));
  AOI211_X1 g442(.A(new_n641_), .B(new_n608_), .C1(new_n626_), .C2(new_n635_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n604_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT72), .B1(new_n622_), .B2(new_n625_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n633_), .A2(new_n634_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n608_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n636_), .A2(new_n642_), .A3(new_n609_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(KEYINPUT13), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G113gat), .B(G141gat), .ZN(new_n652_));
  INV_X1    g451(.A(G197gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT83), .B(G169gat), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n654_), .B(new_n655_), .Z(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n520_), .A2(new_n587_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT82), .ZN(new_n659_));
  INV_X1    g458(.A(new_n587_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(G229gat), .A2(G233gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n466_), .A2(new_n660_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n659_), .A2(new_n665_), .A3(new_n663_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n657_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n666_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n668_), .B(new_n656_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n669_), .A3(KEYINPUT84), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT84), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n671_), .B(new_n657_), .C1(new_n664_), .C2(new_n666_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n645_), .A2(new_n651_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n603_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n265_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n677_), .A2(G1gat), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT38), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n675_), .A2(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n645_), .A2(new_n651_), .A3(KEYINPUT107), .A4(new_n674_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n548_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n454_), .A2(new_n602_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G1gat), .B1(new_n691_), .B2(new_n678_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n680_), .A2(KEYINPUT106), .A3(new_n681_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n679_), .B2(KEYINPUT38), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n682_), .B(new_n692_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1324gat));
  INV_X1    g497(.A(new_n677_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n436_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n583_), .A3(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n690_), .A2(new_n684_), .A3(new_n700_), .A4(new_n685_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT109), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT39), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(G8gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G8gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n701_), .B(new_n708_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1325gat));
  OAI21_X1  g511(.A(G15gat), .B1(new_n691_), .B2(new_n389_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT41), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n677_), .A2(G15gat), .A3(new_n389_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1326gat));
  XNOR2_X1  g515(.A(new_n452_), .B(KEYINPUT111), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n687_), .A2(new_n690_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G22gat), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT42), .ZN(new_n720_));
  INV_X1    g519(.A(G22gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n699_), .A2(new_n721_), .A3(new_n717_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1327gat));
  INV_X1    g522(.A(new_n602_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n454_), .A2(new_n724_), .A3(new_n688_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n676_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(G29gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n265_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT113), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n552_), .A2(new_n557_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n454_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n386_), .A2(new_n392_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n678_), .A3(new_n436_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n451_), .A2(new_n453_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(KEYINPUT43), .A3(new_n558_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n734_), .A2(new_n739_), .A3(new_n602_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n686_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT44), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n265_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n740_), .B2(new_n686_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(KEYINPUT112), .B(new_n744_), .C1(new_n740_), .C2(new_n686_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n731_), .B1(new_n749_), .B2(new_n728_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT114), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n731_), .C1(new_n749_), .C2(new_n728_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1328gat));
  XOR2_X1   g553(.A(KEYINPUT116), .B(KEYINPUT46), .Z(new_n755_));
  INV_X1    g554(.A(G36gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n747_), .A2(new_n748_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n436_), .B1(new_n741_), .B2(KEYINPUT44), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n726_), .A2(G36gat), .A3(new_n436_), .ZN(new_n760_));
  XOR2_X1   g559(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n755_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n759_), .A2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT46), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT117), .B(new_n755_), .C1(new_n759_), .C2(new_n762_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n767_), .A3(new_n768_), .ZN(G1329gat));
  NAND4_X1  g568(.A1(new_n757_), .A2(G43gat), .A3(new_n381_), .A4(new_n742_), .ZN(new_n770_));
  INV_X1    g569(.A(G43gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n726_), .B2(new_n389_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g573(.A(G50gat), .B1(new_n727_), .B2(new_n717_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n452_), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n302_), .B(new_n776_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n777_), .B2(new_n742_), .ZN(G1331gat));
  AND2_X1   g577(.A1(new_n645_), .A2(new_n651_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(new_n674_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n690_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G57gat), .B1(new_n781_), .B2(new_n678_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n780_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n603_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n678_), .A2(G57gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT118), .Z(G1332gat));
  OAI21_X1  g588(.A(G64gat), .B1(new_n781_), .B2(new_n436_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT48), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n436_), .A2(G64gat), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT119), .Z(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n786_), .B2(new_n793_), .ZN(G1333gat));
  OAI21_X1  g593(.A(G71gat), .B1(new_n781_), .B2(new_n389_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT49), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n785_), .A2(new_n566_), .A3(new_n381_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1334gat));
  NAND3_X1  g597(.A1(new_n780_), .A2(new_n690_), .A3(new_n717_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G78gat), .ZN(new_n800_));
  XOR2_X1   g599(.A(KEYINPUT120), .B(KEYINPUT50), .Z(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n785_), .A2(new_n567_), .A3(new_n717_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1335gat));
  AND2_X1   g603(.A1(new_n780_), .A2(new_n725_), .ZN(new_n805_));
  AOI21_X1  g604(.A(G85gat), .B1(new_n805_), .B2(new_n265_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n783_), .A2(new_n740_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n265_), .A2(G85gat), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT121), .Z(new_n810_));
  AOI21_X1  g609(.A(new_n806_), .B1(new_n808_), .B2(new_n810_), .ZN(G1336gat));
  AOI21_X1  g610(.A(G92gat), .B1(new_n805_), .B2(new_n700_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n436_), .A2(new_n489_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n808_), .B2(new_n813_), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n807_), .B2(new_n389_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n805_), .B(new_n381_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(KEYINPUT122), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n817_), .B(new_n819_), .ZN(G1338gat));
  OAI21_X1  g619(.A(G106gat), .B1(new_n807_), .B2(new_n776_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n822_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n805_), .A2(new_n470_), .A3(new_n452_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT123), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n824_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT53), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n823_), .A2(new_n829_), .A3(new_n826_), .A4(new_n824_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1339gat));
  NAND4_X1  g630(.A1(new_n779_), .A2(new_n673_), .A3(new_n724_), .A4(new_n733_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT55), .B1(new_n626_), .B2(new_n635_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n628_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n624_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n633_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n608_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT56), .ZN(new_n841_));
  INV_X1    g640(.A(new_n669_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n663_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n657_), .B1(new_n662_), .B2(new_n843_), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(KEYINPUT125), .Z(new_n845_));
  NAND3_X1  g644(.A1(new_n659_), .A2(new_n665_), .A3(new_n843_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n842_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n848_), .B(new_n608_), .C1(new_n835_), .C2(new_n839_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n841_), .A2(new_n847_), .A3(new_n650_), .A4(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n851_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n558_), .A3(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n841_), .A2(new_n650_), .A3(new_n674_), .A4(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n847_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n688_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(KEYINPUT126), .A2(KEYINPUT57), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n857_), .B(new_n688_), .C1(KEYINPUT126), .C2(KEYINPUT57), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n854_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n834_), .B1(new_n862_), .B2(new_n602_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n700_), .A2(new_n678_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n386_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n863_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867_), .B2(new_n674_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n862_), .A2(new_n602_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n834_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n871_), .A2(KEYINPUT59), .A3(new_n865_), .A4(new_n864_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n673_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n868_), .B1(new_n875_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n779_), .B2(G120gat), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n867_), .B(new_n878_), .C1(new_n877_), .C2(G120gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n779_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n239_), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n867_), .B2(new_n724_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n602_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g683(.A(G134gat), .B1(new_n867_), .B2(new_n689_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n733_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g686(.A(new_n392_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n864_), .A2(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT127), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n863_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n674_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g692(.A(new_n779_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n724_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  AOI21_X1  g698(.A(G162gat), .B1(new_n891_), .B2(new_n689_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n733_), .A2(new_n541_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n891_), .B2(new_n901_), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n436_), .A2(new_n265_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n381_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n717_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n330_), .B1(new_n907_), .B2(new_n674_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n343_), .ZN(new_n909_));
  NOR4_X1   g708(.A1(new_n863_), .A2(new_n673_), .A3(new_n909_), .A4(new_n906_), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT62), .B1(new_n908_), .B2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n863_), .A2(new_n673_), .A3(new_n906_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n330_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n914_), .ZN(G1348gat));
  AOI21_X1  g714(.A(G176gat), .B1(new_n907_), .B2(new_n894_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n863_), .A2(new_n452_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n779_), .A2(new_n331_), .A3(new_n904_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(G1349gat));
  NAND4_X1  g718(.A1(new_n917_), .A2(new_n724_), .A3(new_n381_), .A4(new_n903_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n602_), .A2(new_n323_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n920_), .A2(new_n320_), .B1(new_n907_), .B2(new_n921_), .ZN(G1350gat));
  INV_X1    g721(.A(new_n907_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G190gat), .B1(new_n923_), .B2(new_n733_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n907_), .A2(new_n689_), .A3(new_n322_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1351gat));
  NAND3_X1  g725(.A1(new_n871_), .A2(new_n888_), .A3(new_n903_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n928_), .A2(new_n653_), .A3(new_n674_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G197gat), .B1(new_n927_), .B2(new_n673_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1352gat));
  INV_X1    g730(.A(G204gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n932_), .B1(new_n927_), .B2(new_n779_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n863_), .A2(new_n392_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n934_), .A2(G204gat), .A3(new_n894_), .A4(new_n903_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n927_), .B2(new_n602_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT63), .B(G211gat), .Z(new_n939_));
  NAND4_X1  g738(.A1(new_n934_), .A2(new_n724_), .A3(new_n903_), .A4(new_n939_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1354gat));
  INV_X1    g740(.A(G218gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n934_), .A2(new_n689_), .A3(new_n903_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n733_), .A2(new_n942_), .ZN(new_n944_));
  AOI22_X1  g743(.A1(new_n942_), .A2(new_n943_), .B1(new_n928_), .B2(new_n944_), .ZN(G1355gat));
endmodule


