//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT25), .B(G183gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n207_), .A2(new_n210_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT22), .B1(new_n211_), .B2(KEYINPUT81), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n212_), .B(new_n218_), .C1(new_n219_), .C2(KEYINPUT81), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n205_), .B(new_n206_), .C1(G183gat), .C2(G190gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n214_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n223_), .B(KEYINPUT30), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT82), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(KEYINPUT82), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G71gat), .B(G99gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(G43gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G15gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n230_), .ZN(new_n231_));
  MUX2_X1   g030(.A(new_n225_), .B(new_n226_), .S(new_n231_), .Z(new_n232_));
  XOR2_X1   g031(.A(G127gat), .B(G134gat), .Z(new_n233_));
  XOR2_X1   g032(.A(G113gat), .B(G120gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT31), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n232_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G1gat), .B(G29gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G85gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT0), .B(G57gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G155gat), .B(G162gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(G141gat), .B2(G148gat), .ZN(new_n245_));
  INV_X1    g044(.A(G141gat), .ZN(new_n246_));
  INV_X1    g045(.A(G148gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(KEYINPUT3), .ZN(new_n248_));
  AND3_X1   g047(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT84), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n245_), .A2(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G141gat), .A2(G148gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n252_), .A2(KEYINPUT84), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n243_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n246_), .A2(new_n247_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n243_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n242_), .B1(new_n256_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n235_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n248_), .A2(new_n245_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n249_), .A2(new_n250_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n255_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n260_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n259_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(KEYINPUT1), .B2(new_n243_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(KEYINPUT85), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n263_), .A2(new_n264_), .A3(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n256_), .A2(new_n262_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT97), .B1(new_n273_), .B2(new_n235_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n263_), .A2(new_n264_), .A3(new_n271_), .A4(KEYINPUT97), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT4), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n272_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n241_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n281_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n241_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n284_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n237_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT19), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  INV_X1    g096(.A(G218gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G211gat), .ZN(new_n299_));
  INV_X1    g098(.A(G211gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G218gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n299_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(G197gat), .A2(G204gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT21), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(KEYINPUT21), .A3(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n305_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT88), .B1(new_n303_), .B2(new_n304_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n300_), .A2(G218gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n298_), .A2(G211gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT87), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT88), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n299_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n311_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT89), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n314_), .A2(new_n320_), .A3(new_n324_), .A4(new_n321_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n313_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n207_), .A2(new_n216_), .A3(new_n215_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT93), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n209_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n209_), .A2(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n208_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n214_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT22), .B(G169gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n333_), .B2(new_n212_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n327_), .A2(new_n331_), .B1(new_n221_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n297_), .B1(new_n326_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n313_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n311_), .B1(new_n305_), .B2(new_n318_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n324_), .B1(new_n338_), .B2(new_n314_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n325_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n337_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT94), .B1(new_n341_), .B2(new_n223_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT94), .ZN(new_n343_));
  INV_X1    g142(.A(new_n223_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n326_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n296_), .B(new_n336_), .C1(new_n342_), .C2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT20), .B1(new_n326_), .B2(new_n335_), .ZN(new_n347_));
  AOI211_X1 g146(.A(new_n313_), .B(new_n223_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n295_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G8gat), .B(G36gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT96), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n346_), .A2(new_n355_), .A3(new_n349_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n346_), .A2(new_n355_), .A3(new_n349_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n355_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(KEYINPUT96), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G78gat), .B(G106gat), .Z(new_n366_));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT86), .Z(new_n368_));
  NAND2_X1  g167(.A1(new_n263_), .A2(new_n271_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n341_), .B(new_n368_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT90), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n368_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n273_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n374_), .B1(new_n326_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n371_), .A2(new_n372_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n366_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n366_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n377_), .A4(new_n373_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G22gat), .B(G50gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n369_), .A2(new_n370_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT28), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n386_), .A2(KEYINPUT28), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n385_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n380_), .A2(new_n383_), .B1(KEYINPUT92), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n380_), .A2(new_n383_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n393_), .B(KEYINPUT92), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT101), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n326_), .A2(new_n335_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n348_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT20), .A4(new_n296_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n337_), .B(new_n335_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT20), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n343_), .B1(new_n326_), .B2(new_n344_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n341_), .A2(KEYINPUT94), .A3(new_n223_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n402_), .B1(new_n407_), .B2(new_n296_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n399_), .B1(new_n408_), .B2(new_n356_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n359_), .A2(KEYINPUT27), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n399_), .A3(new_n356_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT102), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n359_), .A2(KEYINPUT27), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n347_), .A2(new_n295_), .A3(new_n348_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n336_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n295_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT101), .B1(new_n417_), .B2(new_n355_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n414_), .A2(new_n418_), .A3(KEYINPUT102), .A4(new_n412_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n365_), .B(new_n398_), .C1(new_n413_), .C2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT103), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n414_), .A2(new_n418_), .A3(new_n412_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT102), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT96), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n350_), .A2(new_n358_), .A3(new_n356_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n426_), .A2(new_n419_), .B1(new_n429_), .B2(new_n364_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(KEYINPUT103), .A3(new_n398_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n293_), .B1(new_n423_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n237_), .B(KEYINPUT83), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n360_), .A2(new_n363_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT99), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n289_), .B2(KEYINPUT98), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n283_), .A2(new_n241_), .A3(new_n285_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n435_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT33), .B1(new_n438_), .B2(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n289_), .A2(KEYINPUT98), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT99), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n280_), .A2(new_n281_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n275_), .A2(new_n276_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n241_), .B1(new_n446_), .B2(new_n282_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n289_), .A2(KEYINPUT33), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  AND4_X1   g247(.A1(new_n434_), .A2(new_n441_), .A3(new_n444_), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT100), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n408_), .A2(KEYINPUT32), .A3(new_n355_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n346_), .A2(new_n349_), .A3(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n291_), .A2(new_n450_), .A3(new_n451_), .A4(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(new_n417_), .B2(new_n452_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT100), .B1(new_n455_), .B2(new_n290_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n398_), .B1(new_n449_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n426_), .A2(new_n419_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n396_), .A2(new_n397_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n394_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n459_), .A2(new_n365_), .A3(new_n290_), .A4(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n433_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n432_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G85gat), .B(G92gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(KEYINPUT8), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT6), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n467_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(KEYINPUT66), .B2(new_n469_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n469_), .A2(KEYINPUT66), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n466_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT67), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT8), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n477_), .A2(new_n478_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n474_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G106gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT10), .B(G99gat), .Z(new_n484_));
  AOI21_X1  g283(.A(new_n470_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n466_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n487_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n482_), .A2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT68), .B(G71gat), .Z(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G78gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT68), .B(G71gat), .ZN(new_n494_));
  INV_X1    g293(.A(G78gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n493_), .B(new_n496_), .C1(KEYINPUT11), .C2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT69), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n498_), .A2(KEYINPUT69), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(KEYINPUT69), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n502_), .A2(KEYINPUT11), .A3(new_n497_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n491_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT12), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n490_), .B(KEYINPUT70), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n482_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n501_), .A2(KEYINPUT12), .A3(new_n504_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n507_), .A2(new_n508_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n482_), .A2(new_n505_), .A3(new_n490_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G230gat), .A2(G233gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT64), .Z(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n515_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n513_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n517_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n514_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n505_), .B1(new_n482_), .B2(new_n490_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G120gat), .B(G148gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(G176gat), .B(G204gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n531_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT13), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(KEYINPUT13), .A3(new_n533_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G29gat), .B(G36gat), .Z(new_n539_));
  XOR2_X1   g338(.A(G43gat), .B(G50gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT15), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543_));
  INV_X1    g342(.A(G1gat), .ZN(new_n544_));
  INV_X1    g343(.A(G8gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G1gat), .B(G8gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n541_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n551_), .B(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n553_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n557_), .A2(KEYINPUT79), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(KEYINPUT79), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n554_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n564_), .A2(KEYINPUT80), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n560_), .B(new_n565_), .Z(new_n566_));
  NOR2_X1   g365(.A1(new_n538_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n465_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n505_), .B(new_n549_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G127gat), .B(G155gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT17), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(KEYINPUT17), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n572_), .A2(new_n578_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(KEYINPUT77), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(KEYINPUT77), .B2(new_n580_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT78), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT34), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n482_), .A2(new_n541_), .A3(new_n490_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n542_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n482_), .B2(new_n509_), .ZN(new_n590_));
  OAI211_X1 g389(.A(KEYINPUT35), .B(new_n587_), .C1(new_n588_), .C2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n510_), .A2(new_n542_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(KEYINPUT35), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n587_), .A2(KEYINPUT35), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n482_), .A2(new_n541_), .A3(new_n490_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n591_), .A2(new_n596_), .A3(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n599_), .B(KEYINPUT36), .Z(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT73), .Z(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n591_), .B2(new_n596_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT37), .B1(new_n601_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n591_), .A2(new_n596_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n602_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n591_), .A2(new_n596_), .A3(new_n600_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n605_), .A2(new_n610_), .A3(KEYINPUT74), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT74), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n613_), .B(KEYINPUT37), .C1(new_n601_), .C2(new_n604_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n611_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n612_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n585_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n569_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT104), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n569_), .A2(KEYINPUT104), .A3(new_n618_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n544_), .A3(new_n291_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT38), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n607_), .A2(new_n609_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n585_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n421_), .A2(new_n422_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT103), .B1(new_n430_), .B2(new_n398_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n292_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n433_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n459_), .A2(new_n365_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n462_), .A2(new_n290_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n454_), .A2(new_n456_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n434_), .A2(new_n441_), .A3(new_n444_), .A4(new_n448_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n462_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n633_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n632_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n629_), .A2(new_n567_), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n290_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n624_), .A2(new_n625_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n626_), .A2(new_n643_), .A3(new_n644_), .ZN(G1324gat));
  XNOR2_X1  g444(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n621_), .A2(new_n545_), .A3(new_n634_), .A4(new_n622_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G8gat), .B1(new_n642_), .B2(new_n430_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n649_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT105), .B(G8gat), .C1(new_n642_), .C2(new_n430_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(KEYINPUT39), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n646_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n656_));
  AND4_X1   g455(.A1(new_n655_), .A2(new_n651_), .A3(new_n647_), .A4(new_n646_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n642_), .B2(new_n633_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT41), .Z(new_n660_));
  INV_X1    g459(.A(G15gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n623_), .A2(new_n661_), .A3(new_n433_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n623_), .A2(new_n664_), .A3(new_n462_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G22gat), .B1(new_n642_), .B2(new_n398_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT42), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1327gat));
  NOR2_X1   g467(.A1(new_n584_), .A2(new_n627_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n569_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G29gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n291_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n585_), .A2(new_n567_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n641_), .B2(new_n617_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n677_), .B(new_n617_), .C1(new_n432_), .C2(new_n464_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT107), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n617_), .B1(new_n432_), .B2(new_n464_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n675_), .B1(new_n685_), .B2(new_n679_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n682_), .A2(new_n683_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n290_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n674_), .B(new_n672_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n688_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT108), .B1(new_n694_), .B2(G29gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n673_), .B1(new_n691_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n430_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n689_), .B2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n430_), .A2(G36gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n670_), .A2(KEYINPUT45), .A3(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT45), .B1(new_n670_), .B2(new_n702_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n697_), .B1(new_n700_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n685_), .A2(new_n679_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n676_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n634_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT44), .B1(new_n681_), .B2(KEYINPUT107), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n688_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT46), .B(new_n705_), .C1(new_n712_), .C2(new_n698_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n707_), .A2(new_n713_), .ZN(G1329gat));
  AOI21_X1  g513(.A(G43gat), .B1(new_n671_), .B2(new_n433_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n237_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G43gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n715_), .B1(new_n689_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(KEYINPUT47), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n721_), .B(new_n715_), .C1(new_n689_), .C2(new_n718_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n671_), .B2(new_n462_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n709_), .A2(G50gat), .A3(new_n462_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n689_), .ZN(G1331gat));
  INV_X1    g525(.A(new_n538_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n566_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n641_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n618_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n291_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n730_), .A2(G57gat), .A3(new_n291_), .A4(new_n629_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n734_), .A2(new_n735_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n733_), .A2(new_n736_), .A3(new_n737_), .ZN(G1332gat));
  NAND2_X1  g537(.A1(new_n730_), .A2(new_n629_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G64gat), .B1(new_n739_), .B2(new_n430_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n430_), .A2(G64gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n731_), .B2(new_n743_), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n739_), .B2(new_n633_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT49), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n633_), .A2(G71gat), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT111), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n731_), .B2(new_n748_), .ZN(G1334gat));
  NAND3_X1  g548(.A1(new_n732_), .A2(new_n495_), .A3(new_n462_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n730_), .A2(new_n462_), .A3(new_n629_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(G78gat), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n751_), .B2(G78gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT112), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n708_), .A2(KEYINPUT114), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n729_), .A2(new_n585_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n685_), .A2(new_n761_), .A3(new_n679_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n758_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n291_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G85gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n641_), .A2(new_n669_), .A3(new_n729_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT113), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n641_), .A2(new_n669_), .A3(new_n729_), .A4(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n290_), .A2(G85gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n765_), .B1(new_n771_), .B2(new_n772_), .ZN(G1336gat));
  AOI21_X1  g572(.A(G92gat), .B1(new_n770_), .B2(new_n634_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n774_), .A2(KEYINPUT115), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(KEYINPUT115), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n634_), .A2(G92gat), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT116), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n775_), .A2(new_n776_), .B1(new_n763_), .B2(new_n778_), .ZN(G1337gat));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n758_), .A2(new_n433_), .A3(new_n760_), .A4(new_n762_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G99gat), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n716_), .A2(new_n484_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n770_), .B2(new_n786_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT117), .B(new_n785_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n780_), .B(KEYINPUT51), .C1(new_n783_), .C2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n780_), .A2(KEYINPUT51), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n782_), .B(new_n791_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1338gat));
  NAND3_X1  g592(.A1(new_n708_), .A2(new_n462_), .A3(new_n760_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(G106gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n794_), .B2(G106gat), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n462_), .A2(new_n483_), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n796_), .A2(new_n797_), .B1(new_n771_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  OAI221_X1 g600(.A(new_n801_), .B1(new_n771_), .B2(new_n798_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  INV_X1    g602(.A(new_n474_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n481_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT8), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n490_), .B(KEYINPUT70), .Z(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n524_), .A2(KEYINPUT12), .B1(new_n810_), .B2(new_n511_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n522_), .B1(new_n811_), .B2(new_n523_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n520_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n813_), .B2(new_n518_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n814_), .B2(KEYINPUT55), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n513_), .B(KEYINPUT55), .C1(new_n520_), .C2(new_n519_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n531_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT56), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n531_), .C1(new_n815_), .C2(new_n817_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n819_), .A2(new_n532_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n550_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n555_), .A2(new_n553_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n564_), .A3(new_n824_), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(KEYINPUT120), .Z(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n564_), .B2(new_n560_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT121), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n822_), .A2(KEYINPUT123), .A3(KEYINPUT58), .A4(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n819_), .A2(new_n532_), .A3(new_n828_), .A4(new_n821_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n829_), .A2(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n835_));
  AOI211_X1 g634(.A(new_n616_), .B(new_n615_), .C1(new_n831_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n819_), .A2(new_n728_), .A3(new_n532_), .A4(new_n821_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n534_), .A2(new_n828_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n840_), .B2(new_n627_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n842_), .B(new_n628_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n585_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n615_), .A2(new_n616_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n536_), .A2(new_n566_), .A3(new_n537_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n584_), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n852_));
  NAND4_X1  g651(.A1(new_n847_), .A2(new_n584_), .A3(new_n848_), .A4(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n846_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n237_), .B1(new_n423_), .B2(new_n431_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n856_), .A2(KEYINPUT59), .A3(new_n291_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n584_), .B1(new_n837_), .B2(new_n844_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n291_), .B(new_n857_), .C1(new_n859_), .C2(new_n854_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n566_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(G113gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n728_), .A2(new_n864_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n863_), .A2(new_n864_), .B1(new_n860_), .B2(new_n865_), .ZN(G1340gat));
  AOI21_X1  g665(.A(new_n727_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n867_));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n727_), .B2(KEYINPUT60), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(KEYINPUT60), .B2(new_n868_), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n867_), .A2(new_n868_), .B1(new_n860_), .B2(new_n870_), .ZN(G1341gat));
  AOI21_X1  g670(.A(new_n585_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n872_));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n584_), .A2(new_n873_), .ZN(new_n874_));
  OAI22_X1  g673(.A1(new_n872_), .A2(new_n873_), .B1(new_n860_), .B2(new_n874_), .ZN(G1342gat));
  AOI21_X1  g674(.A(new_n847_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n876_));
  INV_X1    g675(.A(G134gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n628_), .A2(new_n877_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n876_), .A2(new_n877_), .B1(new_n860_), .B2(new_n878_), .ZN(G1343gat));
  NOR3_X1   g678(.A1(new_n433_), .A2(new_n634_), .A3(new_n398_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n856_), .A2(new_n291_), .A3(new_n880_), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n881_), .A2(G141gat), .A3(new_n566_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G141gat), .B1(new_n881_), .B2(new_n566_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1344gat));
  OR3_X1    g683(.A1(new_n881_), .A2(G148gat), .A3(new_n727_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G148gat), .B1(new_n881_), .B2(new_n727_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1345gat));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  OR3_X1    g687(.A1(new_n881_), .A2(new_n585_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n881_), .B2(new_n585_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1346gat));
  OAI21_X1  g690(.A(G162gat), .B1(new_n881_), .B2(new_n847_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n627_), .A2(G162gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n881_), .B2(new_n893_), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n633_), .A2(new_n291_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n634_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n398_), .B(new_n897_), .C1(new_n859_), .C2(new_n854_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G169gat), .B1(new_n898_), .B2(new_n566_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n898_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n902_), .A2(new_n728_), .A3(new_n333_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT62), .B(G169gat), .C1(new_n898_), .C2(new_n566_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n901_), .A2(new_n903_), .A3(new_n904_), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n902_), .B2(new_n538_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n854_), .B1(new_n845_), .B2(new_n585_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n462_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT124), .B(new_n398_), .C1(new_n859_), .C2(new_n854_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n896_), .A2(new_n212_), .A3(new_n727_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n909_), .A2(KEYINPUT125), .A3(new_n910_), .A4(new_n911_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n906_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NOR3_X1   g715(.A1(new_n898_), .A2(new_n208_), .A3(new_n585_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n909_), .A2(new_n584_), .A3(new_n897_), .A4(new_n910_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n203_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n898_), .B2(new_n847_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n628_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n898_), .B2(new_n921_), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n433_), .A2(new_n635_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n634_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n856_), .A2(new_n728_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(G197gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT126), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n927_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n908_), .A2(new_n924_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n930_), .A2(new_n931_), .A3(G197gat), .A4(new_n728_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n928_), .A2(new_n929_), .A3(new_n932_), .ZN(G1352gat));
  XNOR2_X1  g732(.A(KEYINPUT127), .B(G204gat), .ZN(new_n934_));
  INV_X1    g733(.A(new_n930_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n727_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n930_), .A2(new_n538_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1353gat));
  XNOR2_X1  g738(.A(KEYINPUT63), .B(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n935_), .A2(new_n585_), .A3(new_n940_), .ZN(new_n941_));
  AOI211_X1 g740(.A(KEYINPUT63), .B(G211gat), .C1(new_n930_), .C2(new_n584_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n935_), .B2(new_n847_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n930_), .A2(new_n298_), .A3(new_n628_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1355gat));
endmodule


