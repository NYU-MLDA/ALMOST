//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  INV_X1    g002(.A(G64gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G57gat), .ZN(new_n205_));
  INV_X1    g004(.A(G57gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G64gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT11), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G71gat), .B(G78gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT69), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211_));
  AND2_X1   g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n214_), .B(new_n215_), .C1(new_n202_), .C2(KEYINPUT11), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n210_), .A2(new_n211_), .A3(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n211_), .B1(new_n210_), .B2(new_n216_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n203_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n221_), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT7), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n228_), .A2(new_n229_), .A3(KEYINPUT68), .A4(KEYINPUT7), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n223_), .A2(new_n227_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G85gat), .B(G92gat), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT8), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n235_), .A2(new_n236_), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n221_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT67), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n227_), .A2(new_n223_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n241_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n240_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n206_), .A2(G64gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n204_), .A2(G57gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n215_), .B1(new_n253_), .B2(new_n214_), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n208_), .A2(KEYINPUT69), .A3(new_n209_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT70), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n203_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n210_), .A2(new_n211_), .A3(new_n216_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n244_), .A2(new_n246_), .ZN(new_n260_));
  INV_X1    g059(.A(G85gat), .ZN(new_n261_));
  INV_X1    g060(.A(G92gat), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT9), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n238_), .B2(KEYINPUT9), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT10), .B(G99gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT65), .B1(new_n266_), .B2(new_n229_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n265_), .A2(new_n268_), .A3(G106gat), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n260_), .B(new_n264_), .C1(new_n267_), .C2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n219_), .A2(new_n249_), .A3(new_n259_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT12), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n249_), .A2(new_n270_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n259_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n257_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G230gat), .A2(G233gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n278_), .B(KEYINPUT64), .Z(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT71), .B1(new_n274_), .B2(new_n275_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n219_), .A2(new_n259_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT12), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n249_), .B2(new_n270_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n277_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n279_), .B1(new_n276_), .B2(new_n271_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G120gat), .B(G148gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(G176gat), .B(G204gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT13), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(KEYINPUT13), .A3(new_n296_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT73), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G197gat), .B(G204gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(G211gat), .B(G218gat), .Z(new_n305_));
  INV_X1    g104(.A(KEYINPUT21), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n307_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(G228gat), .A2(G233gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT89), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT2), .ZN(new_n316_));
  INV_X1    g115(.A(G141gat), .ZN(new_n317_));
  INV_X1    g116(.A(G148gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT3), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT2), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(KEYINPUT89), .A3(new_n321_), .ZN(new_n322_));
  OR3_X1    g121(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n316_), .A2(new_n320_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  OR3_X1    g123(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(KEYINPUT1), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n326_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n314_), .B(new_n319_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n328_), .A2(KEYINPUT90), .A3(new_n331_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT29), .A3(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n328_), .A2(new_n331_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n310_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n313_), .A2(new_n336_), .B1(new_n339_), .B2(new_n312_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT91), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n334_), .A2(new_n335_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n338_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT28), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n347_), .A3(new_n338_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G22gat), .B(G50gat), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n350_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n343_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n340_), .B(new_n341_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n346_), .A2(new_n348_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n349_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n340_), .B(new_n342_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n343_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G183gat), .A3(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT84), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n366_), .B2(new_n363_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT81), .B(G183gat), .ZN(new_n368_));
  INV_X1    g167(.A(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(G176gat), .B1(KEYINPUT85), .B2(KEYINPUT22), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G169gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(KEYINPUT25), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT26), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(G190gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(KEYINPUT83), .B2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n380_));
  NOR2_X1   g179(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n381_));
  OAI21_X1  g180(.A(G183gat), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n378_), .A2(KEYINPUT83), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n375_), .A2(new_n379_), .A3(new_n382_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n365_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n363_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT24), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  MUX2_X1   g190(.A(new_n390_), .B(KEYINPUT24), .S(new_n391_), .Z(new_n392_));
  NAND4_X1  g191(.A1(new_n384_), .A2(new_n387_), .A3(new_n388_), .A4(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n374_), .A2(new_n393_), .A3(KEYINPUT30), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G15gat), .B(G43gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n399_), .B(KEYINPUT86), .Z(new_n400_));
  XNOR2_X1  g199(.A(new_n398_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT30), .B1(new_n374_), .B2(new_n393_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n395_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n374_), .A2(new_n393_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n401_), .B1(new_n407_), .B2(new_n394_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n362_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G127gat), .B(G134gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G113gat), .B(G120gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT31), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n402_), .B1(new_n395_), .B2(new_n403_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n401_), .A3(new_n394_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(KEYINPUT87), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n415_), .A2(new_n416_), .A3(KEYINPUT87), .A4(new_n413_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n355_), .A2(new_n361_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n412_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n334_), .A2(new_n422_), .A3(new_n335_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT93), .B1(new_n332_), .B2(new_n422_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT93), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n337_), .A2(new_n426_), .A3(new_n412_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .A4(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT95), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n423_), .A2(KEYINPUT4), .A3(new_n425_), .A4(new_n427_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n424_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n430_), .B(new_n431_), .C1(KEYINPUT4), .C2(new_n423_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G1gat), .B(G29gat), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT0), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT94), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G57gat), .B(G85gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n429_), .A2(new_n432_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT19), .ZN(new_n444_));
  OR2_X1    g243(.A1(G183gat), .A2(G190gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n387_), .A2(new_n388_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT92), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n387_), .A2(new_n448_), .A3(new_n388_), .A4(new_n445_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G169gat), .ZN(new_n450_));
  INV_X1    g249(.A(G176gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n447_), .A2(new_n449_), .A3(new_n389_), .A4(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT25), .B(G183gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n377_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n378_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n367_), .A2(new_n392_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n311_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT20), .B1(new_n405_), .B2(new_n310_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n444_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n453_), .A2(new_n457_), .A3(new_n311_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n405_), .A2(new_n310_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n444_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT20), .A4(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT18), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n460_), .A2(new_n471_), .A3(new_n464_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n423_), .A2(new_n431_), .A3(new_n425_), .A4(new_n427_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n438_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n423_), .A2(KEYINPUT4), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(new_n431_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n477_), .B2(new_n430_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n429_), .A2(KEYINPUT33), .A3(new_n432_), .A4(new_n439_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n442_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n463_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT20), .A4(new_n444_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n471_), .A2(KEYINPUT32), .ZN(new_n485_));
  MUX2_X1   g284(.A(new_n484_), .B(new_n465_), .S(new_n485_), .Z(new_n486_));
  INV_X1    g285(.A(new_n440_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n439_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n421_), .B1(new_n481_), .B2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n487_), .A2(new_n488_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n353_), .A2(new_n354_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n360_), .B1(new_n359_), .B2(new_n343_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n420_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n418_), .A2(new_n419_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n355_), .A2(new_n361_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n491_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n473_), .A2(KEYINPUT27), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT96), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n472_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n460_), .A2(new_n464_), .A3(KEYINPUT96), .A4(new_n471_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n482_), .A2(new_n469_), .A3(new_n483_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT27), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n490_), .B1(new_n497_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT15), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT76), .B(G8gat), .ZN(new_n511_));
  INV_X1    g310(.A(G1gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n514_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n515_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n510_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n509_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT77), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n521_), .A2(new_n526_), .A3(new_n509_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n521_), .A2(new_n509_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT77), .B1(new_n521_), .B2(new_n509_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n525_), .B(KEYINPUT80), .C1(new_n530_), .C2(new_n524_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT78), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n533_), .B(KEYINPUT79), .Z(new_n534_));
  XNOR2_X1  g333(.A(G169gat), .B(G197gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n531_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT37), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT35), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n273_), .B2(new_n510_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n249_), .A2(new_n270_), .A3(new_n509_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(KEYINPUT35), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT74), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT74), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n543_), .A2(KEYINPUT74), .A3(new_n544_), .A4(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT75), .ZN(new_n554_));
  XOR2_X1   g353(.A(G134gat), .B(G162gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT36), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n556_), .B(KEYINPUT36), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n552_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n539_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n558_), .B(KEYINPUT37), .C1(new_n552_), .C2(new_n561_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n280_), .A2(new_n282_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n521_), .B(new_n567_), .Z(new_n568_));
  AND2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT16), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n569_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n568_), .B2(new_n566_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n274_), .A2(new_n275_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(new_n568_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n568_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n574_), .B(KEYINPUT17), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n565_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR4_X1   g384(.A1(new_n303_), .A2(new_n506_), .A3(new_n538_), .A4(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n512_), .A3(new_n491_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT38), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n481_), .A2(new_n489_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n421_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n487_), .A2(new_n488_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n355_), .A2(new_n361_), .A3(new_n495_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n495_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n592_), .B(new_n505_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n301_), .A2(new_n538_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n559_), .A2(new_n562_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n583_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n512_), .B1(new_n601_), .B2(new_n491_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT97), .Z(new_n603_));
  NAND2_X1  g402(.A1(new_n588_), .A2(new_n603_), .ZN(G1324gat));
  INV_X1    g403(.A(new_n505_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n586_), .A2(new_n511_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT98), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(new_n605_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(G8gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT39), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(KEYINPUT39), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g412(.A1(new_n601_), .A2(new_n495_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G15gat), .ZN(new_n615_));
  XOR2_X1   g414(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n586_), .A2(new_n619_), .A3(new_n495_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT100), .Z(G1326gat));
  INV_X1    g421(.A(G22gat), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n492_), .A2(new_n493_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n601_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n586_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1327gat));
  NAND2_X1  g429(.A1(new_n583_), .A2(new_n599_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT106), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n598_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n491_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  INV_X1    g435(.A(new_n565_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n638_), .B2(KEYINPUT102), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n640_), .B(KEYINPUT43), .C1(new_n506_), .C2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n642_), .A2(KEYINPUT44), .A3(new_n583_), .A4(new_n597_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n583_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n647_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n597_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n649_), .A2(G29gat), .A3(new_n491_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n596_), .A2(new_n565_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT43), .B1(new_n651_), .B2(new_n640_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n638_), .A2(KEYINPUT102), .A3(new_n636_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n583_), .B(new_n597_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT103), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n647_), .A2(new_n656_), .A3(new_n597_), .ZN(new_n657_));
  XOR2_X1   g456(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n635_), .B1(new_n650_), .B2(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n634_), .A2(new_n663_), .A3(new_n605_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n665_));
  AOI21_X1  g464(.A(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n649_), .A2(new_n659_), .A3(KEYINPUT107), .A4(new_n605_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n662_), .A2(new_n663_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n658_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n654_), .B2(KEYINPUT103), .ZN(new_n672_));
  AOI22_X1  g471(.A1(new_n657_), .A2(new_n672_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT107), .B1(new_n673_), .B2(new_n605_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n661_), .B(new_n667_), .C1(new_n670_), .C2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n649_), .A2(new_n659_), .A3(new_n605_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n661_), .B1(new_n680_), .B2(new_n667_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n676_), .A2(new_n681_), .ZN(G1329gat));
  NAND3_X1  g481(.A1(new_n673_), .A2(G43gat), .A3(new_n495_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n633_), .A2(new_n420_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(G43gat), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g485(.A(G50gat), .B1(new_n634_), .B2(new_n625_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n649_), .A2(G50gat), .A3(new_n625_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n659_), .ZN(G1331gat));
  INV_X1    g488(.A(new_n301_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n537_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(new_n596_), .A3(new_n584_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G57gat), .B1(new_n692_), .B2(new_n491_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT110), .Z(new_n694_));
  NOR3_X1   g493(.A1(new_n302_), .A2(new_n506_), .A3(new_n537_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(new_n600_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(KEYINPUT111), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(KEYINPUT111), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n592_), .A2(new_n206_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n694_), .B1(new_n700_), .B2(new_n701_), .ZN(G1332gat));
  NAND3_X1  g501(.A1(new_n692_), .A2(new_n204_), .A3(new_n605_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n605_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G64gat), .ZN(new_n706_));
  AOI211_X1 g505(.A(KEYINPUT48), .B(new_n204_), .C1(new_n700_), .C2(new_n605_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(G1333gat));
  OAI21_X1  g507(.A(G71gat), .B1(new_n699_), .B2(new_n420_), .ZN(new_n709_));
  XOR2_X1   g508(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n710_));
  OR2_X1    g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  INV_X1    g511(.A(G71gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n692_), .A2(new_n713_), .A3(new_n495_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n712_), .A3(new_n714_), .ZN(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n692_), .A2(new_n716_), .A3(new_n625_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n700_), .A2(new_n625_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G78gat), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT50), .B(new_n716_), .C1(new_n700_), .C2(new_n625_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1335gat));
  AND2_X1   g521(.A1(new_n647_), .A2(new_n691_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n592_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n695_), .A2(new_n632_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n261_), .A3(new_n491_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1336gat));
  OAI21_X1  g527(.A(G92gat), .B1(new_n724_), .B2(new_n505_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n262_), .A3(new_n605_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1337gat));
  NOR2_X1   g530(.A1(new_n420_), .A2(new_n265_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT114), .B1(new_n726_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n723_), .A2(new_n495_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n734_), .A2(KEYINPUT113), .A3(G99gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT113), .B1(new_n734_), .B2(G99gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n733_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g537(.A1(new_n726_), .A2(new_n229_), .A3(new_n625_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n723_), .A2(new_n625_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(G106gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT52), .B(new_n229_), .C1(new_n723_), .C2(new_n625_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g544(.A(KEYINPUT125), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n605_), .A2(new_n592_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n593_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT123), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT59), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n536_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n530_), .A2(new_n524_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n752_), .B(new_n753_), .C1(new_n524_), .C2(new_n523_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n530_), .A2(new_n524_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n524_), .B2(new_n523_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n756_), .B2(new_n752_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT119), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT119), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n754_), .B(new_n759_), .C1(new_n756_), .C2(new_n752_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n294_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT120), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n758_), .A2(new_n294_), .A3(KEYINPUT120), .A4(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n279_), .B1(new_n277_), .B2(new_n285_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n286_), .B2(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n277_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n770_));
  AND3_X1   g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n295_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n295_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(KEYINPUT121), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n777_), .B(KEYINPUT56), .C1(new_n773_), .C2(new_n295_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT58), .B(new_n765_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT122), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n765_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n768_), .A2(new_n770_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT117), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n293_), .B1(new_n788_), .B2(new_n767_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n777_), .B1(new_n789_), .B2(KEYINPUT56), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n773_), .A2(new_n295_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT121), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n793_), .A3(new_n774_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(KEYINPUT122), .A3(KEYINPUT58), .A4(new_n765_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n781_), .A2(new_n784_), .A3(new_n565_), .A4(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n797_));
  NOR2_X1   g596(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n789_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n294_), .A2(new_n537_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n294_), .A2(KEYINPUT115), .A3(new_n537_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n797_), .A2(new_n799_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n297_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n599_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n796_), .A2(KEYINPUT124), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n806_), .A2(KEYINPUT57), .A3(new_n807_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT124), .B1(new_n796_), .B2(new_n810_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n583_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n690_), .A2(new_n538_), .A3(new_n584_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n816_), .A2(KEYINPUT54), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(KEYINPUT54), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n751_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n819_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n796_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n583_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT59), .B1(new_n823_), .B2(new_n748_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n746_), .B1(new_n820_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n796_), .A2(new_n810_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n812_), .A3(new_n811_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n821_), .B1(new_n830_), .B2(new_n583_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT125), .B(new_n824_), .C1(new_n831_), .C2(new_n751_), .ZN(new_n832_));
  INV_X1    g631(.A(G113gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n538_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n826_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n823_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n748_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n838_), .B2(new_n538_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n835_), .A2(new_n839_), .ZN(G1340gat));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n841_));
  INV_X1    g640(.A(G120gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n301_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n836_), .A2(new_n837_), .A3(new_n844_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n820_), .A2(new_n825_), .A3(new_n302_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n842_), .ZN(G1341gat));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n583_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n826_), .A2(new_n832_), .A3(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n838_), .B2(new_n583_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n637_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n826_), .A2(new_n832_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n838_), .B2(new_n807_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n823_), .A2(new_n494_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n747_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n538_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n317_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n302_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n318_), .ZN(G1345gat));
  NOR2_X1   g662(.A1(new_n859_), .A2(new_n583_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G155gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  OAI21_X1  g665(.A(G162gat), .B1(new_n859_), .B2(new_n637_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n807_), .A2(G162gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n859_), .B2(new_n868_), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n815_), .A2(new_n819_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n505_), .A2(new_n491_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n495_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n625_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n870_), .A2(new_n450_), .A3(new_n537_), .A4(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n870_), .A2(new_n537_), .A3(new_n873_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n875_), .A2(new_n876_), .A3(G169gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n875_), .B2(G169gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n874_), .B1(new_n877_), .B2(new_n878_), .ZN(G1348gat));
  NAND3_X1  g678(.A1(new_n870_), .A2(new_n301_), .A3(new_n873_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n823_), .A2(new_n625_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n302_), .A2(new_n451_), .A3(new_n872_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n880_), .A2(new_n451_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  NAND2_X1  g682(.A1(new_n870_), .A2(new_n873_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n884_), .A2(new_n583_), .A3(new_n454_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n881_), .A2(new_n646_), .A3(new_n495_), .A4(new_n871_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n368_), .B2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n884_), .B2(new_n637_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n599_), .A2(new_n378_), .A3(new_n455_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n884_), .B2(new_n889_), .ZN(G1351gat));
  AND2_X1   g689(.A1(new_n858_), .A2(new_n871_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n537_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n303_), .ZN(new_n894_));
  INV_X1    g693(.A(G204gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(KEYINPUT126), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n894_), .B(new_n896_), .ZN(G1353gat));
  AOI21_X1  g696(.A(new_n583_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT127), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n891_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n900_), .B(new_n902_), .ZN(G1354gat));
  INV_X1    g702(.A(G218gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n891_), .A2(new_n904_), .A3(new_n599_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n891_), .A2(new_n565_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n904_), .ZN(G1355gat));
endmodule


