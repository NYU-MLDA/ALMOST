//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_;
  XNOR2_X1  g000(.A(G1gat), .B(G8gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT71), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G1gat), .A2(G8gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT14), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n202_), .A2(KEYINPUT71), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n202_), .A2(KEYINPUT71), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n209_), .A2(new_n206_), .A3(new_n204_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n212_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT74), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n212_), .A2(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n215_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT74), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n215_), .B(new_n225_), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n226_), .A2(KEYINPUT75), .A3(new_n212_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT75), .B1(new_n226_), .B2(new_n212_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n224_), .B1(new_n212_), .B2(new_n215_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n222_), .A2(new_n224_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G113gat), .B(G141gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G169gat), .B(G197gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n232_), .B(new_n233_), .Z(new_n234_));
  XOR2_X1   g033(.A(new_n231_), .B(new_n234_), .Z(new_n235_));
  XNOR2_X1  g034(.A(G8gat), .B(G36gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT18), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G64gat), .B(G92gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G169gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT95), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n243_), .B2(G176gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT96), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G183gat), .A2(G190gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT23), .ZN(new_n248_));
  OR2_X1    g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n244_), .A2(new_n245_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT25), .B(G183gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G169gat), .ZN(new_n255_));
  INV_X1    g054(.A(G176gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT24), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT24), .A3(new_n241_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n254_), .A2(new_n248_), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n251_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G197gat), .B(G204gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G211gat), .B(G218gat), .Z(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT21), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G204gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n268_));
  OAI211_X1 g067(.A(KEYINPUT21), .B(new_n268_), .C1(new_n263_), .C2(KEYINPUT88), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n264_), .B1(new_n262_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT90), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(KEYINPUT90), .A3(new_n271_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n266_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n261_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT19), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT20), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT76), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT22), .B1(new_n283_), .B2(new_n255_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT22), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(KEYINPUT76), .A3(G169gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n256_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT77), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n248_), .A2(new_n249_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n241_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n260_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n282_), .B1(new_n292_), .B2(new_n276_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n278_), .A2(new_n281_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT101), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n278_), .A2(KEYINPUT101), .A3(new_n281_), .A4(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n261_), .A2(KEYINPUT100), .ZN(new_n299_));
  INV_X1    g098(.A(new_n260_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n246_), .B2(new_n250_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT100), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n276_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n282_), .B1(new_n277_), .B2(new_n291_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n281_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n240_), .B1(new_n298_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n301_), .A2(new_n276_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT20), .B1(new_n277_), .B2(new_n291_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n280_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n301_), .A2(new_n276_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n305_), .A3(new_n281_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n312_), .A3(new_n239_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(KEYINPUT27), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(KEYINPUT1), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT83), .ZN(new_n318_));
  INV_X1    g117(.A(G155gat), .ZN(new_n319_));
  INV_X1    g118(.A(G162gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n321_), .A2(new_n322_), .B1(KEYINPUT1), .B2(new_n316_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT84), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n317_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n324_), .B2(new_n323_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT82), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n321_), .A2(new_n322_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n327_), .B(KEYINPUT3), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n329_), .B(KEYINPUT2), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n332_), .B(new_n316_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n331_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G127gat), .B(G134gat), .Z(new_n340_));
  XOR2_X1   g139(.A(G113gat), .B(G120gat), .Z(new_n341_));
  XOR2_X1   g140(.A(new_n340_), .B(new_n341_), .Z(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n343_), .A2(KEYINPUT4), .ZN(new_n344_));
  INV_X1    g143(.A(new_n342_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n331_), .A2(new_n338_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(KEYINPUT4), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n315_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n346_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n349_), .A2(new_n315_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G85gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT0), .B(G57gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  OR3_X1    g153(.A1(new_n348_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT97), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n313_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT97), .A4(new_n239_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n310_), .A2(new_n312_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n240_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n314_), .A2(new_n358_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n368_), .B(KEYINPUT87), .Z(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n331_), .B2(new_n338_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n277_), .B(new_n370_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n373_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT91), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n372_), .A2(new_n373_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n276_), .A2(new_n369_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT91), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .A4(new_n375_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n368_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(new_n372_), .B2(new_n276_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(KEYINPUT92), .B(new_n383_), .C1(new_n372_), .C2(new_n276_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT93), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n331_), .A2(new_n338_), .A3(new_n371_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT28), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G22gat), .B(G50gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n394_), .B(new_n395_), .Z(new_n396_));
  AOI22_X1  g195(.A1(new_n377_), .A2(new_n381_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n391_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT93), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n382_), .A2(new_n398_), .A3(new_n388_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n392_), .B(new_n396_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n391_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n396_), .B1(new_n397_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n389_), .A2(new_n402_), .A3(new_n391_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407_));
  INV_X1    g206(.A(G43gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n291_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT30), .ZN(new_n414_));
  INV_X1    g213(.A(new_n409_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n290_), .A2(new_n415_), .A3(new_n260_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n410_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n414_), .B1(new_n410_), .B2(new_n416_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT78), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n342_), .B(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n423_), .B2(KEYINPUT80), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n419_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(KEYINPUT78), .A3(new_n417_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n428_), .A2(KEYINPUT80), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n426_), .B(KEYINPUT81), .C1(new_n429_), .C2(new_n423_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT81), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n423_), .B1(new_n428_), .B2(KEYINPUT80), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n425_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n401_), .A2(new_n406_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n401_), .B2(new_n406_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n367_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n401_), .A2(new_n406_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n239_), .A2(KEYINPUT32), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n310_), .A2(new_n312_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT99), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n440_), .A2(new_n441_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n357_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n298_), .A2(new_n306_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(new_n439_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT98), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(KEYINPUT33), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n356_), .B(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n344_), .A2(new_n315_), .A3(new_n347_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n354_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n450_), .B(new_n451_), .C1(new_n315_), .C2(new_n349_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n360_), .A2(new_n363_), .A3(new_n361_), .A4(new_n452_), .ZN(new_n453_));
  OAI22_X1  g252(.A1(new_n444_), .A2(new_n446_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n434_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n438_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n235_), .B1(new_n437_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G85gat), .ZN(new_n458_));
  INV_X1    g257(.A(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT9), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n471_));
  INV_X1    g270(.A(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n464_), .A2(new_n465_), .A3(new_n470_), .A4(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(KEYINPUT8), .B(new_n462_), .C1(new_n479_), .C2(new_n470_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n482_));
  INV_X1    g281(.A(G99gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n483_), .A3(new_n472_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n468_), .B1(G99gat), .B2(G106gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n476_), .B(new_n484_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n481_), .B1(new_n487_), .B2(new_n463_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n475_), .B1(new_n480_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT64), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(new_n475_), .C1(new_n480_), .C2(new_n488_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n215_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G232gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT34), .ZN(new_n495_));
  INV_X1    g294(.A(new_n489_), .ZN(new_n496_));
  OAI221_X1 g295(.A(new_n493_), .B1(KEYINPUT35), .B2(new_n495_), .C1(new_n226_), .C2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n495_), .A2(KEYINPUT35), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n497_), .A2(new_n498_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G190gat), .B(G218gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(G134gat), .B(G162gat), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n503_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT36), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT69), .Z(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n504_), .A2(KEYINPUT36), .A3(new_n505_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(new_n506_), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n510_), .B(KEYINPUT70), .Z(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT37), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n510_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n212_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G71gat), .B(G78gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n525_));
  INV_X1    g324(.A(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT67), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n531_), .B(new_n524_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n521_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G127gat), .B(G155gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT16), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n520_), .A2(new_n532_), .A3(new_n530_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT72), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n521_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n529_), .A2(KEYINPUT65), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT65), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(new_n524_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n520_), .A2(KEYINPUT72), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n538_), .B(KEYINPUT17), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n549_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n542_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT73), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n518_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n490_), .A2(new_n492_), .A3(new_n548_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n548_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n490_), .A2(new_n492_), .A3(new_n548_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n533_), .A2(KEYINPUT12), .A3(new_n489_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n563_), .B(new_n564_), .C1(new_n561_), .C2(KEYINPUT12), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n562_), .B(KEYINPUT66), .C1(new_n565_), .C2(new_n559_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT66), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n567_), .B(new_n559_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT5), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(KEYINPUT68), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n566_), .B(new_n568_), .C1(KEYINPUT68), .C2(new_n574_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT13), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(KEYINPUT13), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n557_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n457_), .A2(new_n581_), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n582_), .A2(G1gat), .A3(new_n358_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT38), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT102), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(new_n579_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n235_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT103), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(new_n555_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n508_), .A2(new_n516_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n437_), .B2(new_n456_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n357_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n598_), .A2(G1gat), .B1(new_n584_), .B2(new_n583_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n586_), .A2(new_n599_), .ZN(G1324gat));
  AND2_X1   g399(.A1(new_n314_), .A2(new_n366_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n582_), .A2(G8gat), .A3(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G8gat), .B1(new_n596_), .B2(new_n601_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT39), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n605_), .B(G8gat), .C1(new_n596_), .C2(new_n601_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n602_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n607_), .B(new_n609_), .ZN(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n596_), .B2(new_n455_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT41), .Z(new_n612_));
  INV_X1    g411(.A(new_n582_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n412_), .A3(new_n434_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(G1326gat));
  OR3_X1    g414(.A1(new_n582_), .A2(G22gat), .A3(new_n438_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n438_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n597_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n619_));
  AND3_X1   g418(.A1(new_n618_), .A2(G22gat), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n618_), .B2(G22gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n616_), .B1(new_n620_), .B2(new_n621_), .ZN(G1327gat));
  INV_X1    g421(.A(new_n556_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n457_), .A2(new_n594_), .A3(new_n623_), .A4(new_n587_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n624_), .A2(G29gat), .A3(new_n358_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n589_), .B(KEYINPUT103), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n437_), .A2(new_n456_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n518_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT43), .B(new_n518_), .C1(new_n437_), .C2(new_n456_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n623_), .B(new_n626_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT107), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT107), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n632_), .A2(new_n636_), .A3(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n632_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n358_), .B1(new_n639_), .B2(KEYINPUT44), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(KEYINPUT108), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G29gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT108), .B1(new_n638_), .B2(new_n640_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n625_), .B1(new_n642_), .B2(new_n643_), .ZN(G1328gat));
  NOR3_X1   g443(.A1(new_n624_), .A2(G36gat), .A3(new_n601_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT45), .Z(new_n646_));
  INV_X1    g445(.A(new_n601_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n632_), .B2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n650_));
  INV_X1    g449(.A(G36gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n646_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT46), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT46), .B(new_n646_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1329gat));
  NAND2_X1  g455(.A1(new_n639_), .A2(KEYINPUT44), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n455_), .A2(new_n408_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n637_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n636_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n657_), .B(new_n658_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n408_), .B1(new_n624_), .B2(new_n455_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT47), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT47), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n665_), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1330gat));
  INV_X1    g466(.A(G50gat), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n438_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n657_), .B(new_n669_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n624_), .B2(new_n438_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT109), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(new_n674_), .A3(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1331gat));
  AOI21_X1  g475(.A(new_n588_), .B1(new_n437_), .B2(new_n456_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n587_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n518_), .A2(new_n677_), .A3(new_n556_), .A4(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G57gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n357_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n587_), .A2(new_n588_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n595_), .A2(new_n556_), .A3(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(new_n357_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n684_), .B2(new_n680_), .ZN(G1332gat));
  INV_X1    g484(.A(G64gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n683_), .B2(new_n647_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT48), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n679_), .A2(new_n686_), .A3(new_n647_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1333gat));
  INV_X1    g489(.A(G71gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n683_), .B2(new_n434_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT49), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n679_), .A2(new_n691_), .A3(new_n434_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1334gat));
  INV_X1    g494(.A(G78gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n683_), .B2(new_n617_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT50), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n679_), .A2(new_n696_), .A3(new_n617_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1335gat));
  INV_X1    g499(.A(new_n630_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n631_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(new_n623_), .A3(new_n682_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G85gat), .B1(new_n704_), .B2(new_n358_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n587_), .A2(new_n593_), .A3(new_n556_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n677_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n458_), .A3(new_n357_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(G1336gat));
  OAI21_X1  g509(.A(G92gat), .B1(new_n704_), .B2(new_n601_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(new_n459_), .A3(new_n647_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT110), .ZN(G1337gat));
  NAND4_X1  g513(.A1(new_n708_), .A2(new_n434_), .A3(new_n471_), .A4(new_n473_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT111), .ZN(new_n716_));
  OAI21_X1  g515(.A(G99gat), .B1(new_n704_), .B2(new_n455_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g518(.A1(new_n708_), .A2(new_n472_), .A3(new_n617_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n703_), .A2(new_n617_), .A3(new_n623_), .A4(new_n682_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(G106gat), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n721_), .B2(G106gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n720_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT53), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n728_), .B(new_n720_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1339gat));
  NAND2_X1  g529(.A1(new_n601_), .A2(new_n357_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n731_), .A2(new_n617_), .A3(new_n455_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT59), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT54), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n581_), .B2(new_n235_), .ZN(new_n736_));
  NOR4_X1   g535(.A1(new_n678_), .A2(new_n557_), .A3(KEYINPUT54), .A4(new_n588_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n565_), .A2(new_n559_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT112), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n565_), .A2(new_n741_), .A3(new_n559_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT55), .B1(new_n565_), .B2(new_n559_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n561_), .A2(KEYINPUT12), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n563_), .A2(new_n564_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .A4(new_n558_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n743_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n574_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n750_), .A2(KEYINPUT113), .A3(new_n752_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n740_), .A2(new_n742_), .B1(new_n744_), .B2(new_n748_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n754_), .B2(new_n574_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  INV_X1    g555(.A(new_n752_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(new_n755_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n569_), .A2(new_n574_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n235_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n222_), .A2(new_n223_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n223_), .B1(new_n212_), .B2(new_n215_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n234_), .B1(new_n229_), .B2(new_n765_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n231_), .A2(new_n234_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n576_), .A2(new_n577_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT114), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n576_), .A2(new_n770_), .A3(new_n577_), .A4(new_n767_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n594_), .B1(new_n763_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n760_), .A2(new_n767_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT56), .B1(new_n750_), .B2(new_n573_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n754_), .A2(new_n757_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n518_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT58), .B(new_n775_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n773_), .A2(KEYINPUT57), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n773_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n769_), .A2(new_n771_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n786_), .A2(KEYINPUT115), .A3(new_n594_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n781_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n623_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n738_), .B1(new_n789_), .B2(KEYINPUT117), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT115), .B1(new_n786_), .B2(new_n594_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n763_), .A2(new_n772_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(new_n783_), .A3(new_n593_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n793_), .A3(new_n782_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n556_), .B1(new_n794_), .B2(new_n781_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n734_), .B1(new_n790_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n738_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n788_), .A2(new_n555_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n733_), .B1(new_n801_), .B2(new_n732_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n798_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n588_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(G113gat), .ZN(new_n805_));
  INV_X1    g604(.A(new_n555_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n794_), .B2(new_n781_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n732_), .B1(new_n807_), .B2(new_n738_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n808_), .A2(G113gat), .A3(new_n235_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n805_), .A2(new_n809_), .ZN(G1340gat));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(KEYINPUT59), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n678_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n813_), .B2(new_n798_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n799_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n789_), .A2(KEYINPUT117), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n733_), .B(new_n732_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(KEYINPUT118), .A3(new_n678_), .A4(new_n812_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(new_n818_), .A3(G120gat), .ZN(new_n819_));
  INV_X1    g618(.A(new_n808_), .ZN(new_n820_));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n820_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n821_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n823_), .ZN(G1341gat));
  AOI21_X1  g623(.A(G127gat), .B1(new_n820_), .B2(new_n556_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n806_), .A2(G127gat), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT119), .Z(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n803_), .B2(new_n827_), .ZN(G1342gat));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  INV_X1    g628(.A(G134gat), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n518_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n798_), .A2(new_n802_), .A3(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n594_), .B(new_n732_), .C1(new_n807_), .C2(new_n738_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n830_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT120), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n837_), .A3(new_n830_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n829_), .B1(new_n833_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n817_), .A2(new_n812_), .A3(new_n831_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n841_), .A2(KEYINPUT121), .A3(new_n836_), .A4(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1343gat));
  NOR2_X1   g642(.A1(new_n807_), .A2(new_n738_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n436_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n731_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT122), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849_));
  NOR4_X1   g648(.A1(new_n844_), .A2(new_n849_), .A3(new_n845_), .A4(new_n731_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n588_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G141gat), .ZN(new_n852_));
  INV_X1    g651(.A(G141gat), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n853_), .B(new_n588_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1344gat));
  OAI21_X1  g654(.A(new_n678_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G148gat), .ZN(new_n857_));
  INV_X1    g656(.A(G148gat), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n858_), .B(new_n678_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1345gat));
  OAI21_X1  g659(.A(new_n556_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n862_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n556_), .B(new_n864_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1346gat));
  OAI211_X1 g665(.A(new_n320_), .B(new_n594_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n846_), .A2(new_n847_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n849_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n850_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n518_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n871_), .B2(new_n320_), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n601_), .A2(new_n357_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n434_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n876_), .A3(new_n434_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n617_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT126), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n883_), .B(new_n880_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n235_), .A2(new_n243_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT127), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n882_), .A2(new_n884_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT124), .B1(new_n878_), .B2(new_n588_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  AOI211_X1 g688(.A(new_n889_), .B(new_n235_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n438_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n797_), .B2(new_n790_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n255_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n892_), .A2(new_n255_), .A3(new_n894_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n887_), .B1(new_n896_), .B2(new_n897_), .ZN(G1348gat));
  NAND3_X1  g697(.A1(new_n882_), .A2(new_n884_), .A3(new_n678_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n844_), .A2(new_n617_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n879_), .A2(new_n256_), .A3(new_n587_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n899_), .A2(new_n256_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  NOR2_X1   g701(.A1(new_n879_), .A2(new_n623_), .ZN(new_n903_));
  AOI21_X1  g702(.A(G183gat), .B1(new_n900_), .B2(new_n903_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n882_), .A2(new_n884_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n555_), .A2(new_n252_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n904_), .B1(new_n905_), .B2(new_n907_), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n882_), .A2(new_n884_), .A3(new_n629_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G190gat), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n882_), .A2(new_n884_), .A3(new_n253_), .A4(new_n594_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1351gat));
  NAND2_X1  g711(.A1(new_n846_), .A2(new_n873_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n235_), .ZN(new_n914_));
  INV_X1    g713(.A(G197gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1352gat));
  NOR2_X1   g715(.A1(new_n913_), .A2(new_n587_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(new_n267_), .ZN(G1353gat));
  INV_X1    g717(.A(new_n913_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT63), .B(G211gat), .Z(new_n920_));
  NAND3_X1  g719(.A1(new_n919_), .A2(new_n806_), .A3(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n922_), .B1(new_n913_), .B2(new_n555_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1354gat));
  OR3_X1    g723(.A1(new_n913_), .A2(G218gat), .A3(new_n593_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G218gat), .B1(new_n913_), .B2(new_n518_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1355gat));
endmodule


