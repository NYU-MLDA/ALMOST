//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G64gat), .ZN(new_n204_));
  INV_X1    g003(.A(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT93), .Z(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT19), .Z(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G197gat), .B(G204gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(G211gat), .B(G218gat), .Z(new_n213_));
  INV_X1    g012(.A(KEYINPUT21), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G211gat), .B(G218gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT21), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n215_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n225_), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n220_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT81), .B(G183gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n220_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT83), .B(G176gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(new_n221_), .B2(KEYINPUT22), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G169gat), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n238_), .B(new_n240_), .C1(new_n241_), .C2(new_n239_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n225_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n244_), .A2(KEYINPUT84), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(KEYINPUT84), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n218_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT96), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT20), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT25), .B(G183gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n228_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n227_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n241_), .A2(new_n238_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n225_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT95), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n255_), .A2(KEYINPUT95), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n253_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n215_), .B(new_n217_), .Z(new_n262_));
  AOI21_X1  g061(.A(new_n250_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n211_), .B1(new_n249_), .B2(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n244_), .A2(KEYINPUT84), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n244_), .A2(KEYINPUT84), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n262_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT94), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT20), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n218_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n267_), .B2(KEYINPUT20), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n271_), .A2(new_n210_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n207_), .B1(new_n264_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT100), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT100), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n276_), .B(new_n207_), .C1(new_n264_), .C2(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n249_), .A2(new_n211_), .A3(new_n263_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n210_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n206_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n281_), .A2(KEYINPUT27), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n280_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n207_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n281_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n278_), .A2(new_n282_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT88), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293_));
  AND2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n293_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT89), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n288_), .B(new_n290_), .C1(new_n295_), .C2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n294_), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n288_), .B(KEYINPUT2), .Z(new_n304_));
  NOR2_X1   g103(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n289_), .B(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n292_), .B(new_n303_), .C1(new_n304_), .C2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n299_), .A2(new_n302_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT97), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT97), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n299_), .A2(new_n310_), .A3(new_n302_), .A4(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n299_), .A2(new_n307_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n300_), .A2(new_n301_), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(new_n302_), .B2(KEYINPUT86), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n309_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT4), .B1(new_n312_), .B2(new_n315_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(new_n317_), .B2(KEYINPUT4), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n318_), .B(KEYINPUT98), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n320_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G1gat), .B(G29gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT0), .ZN(new_n327_));
  INV_X1    g126(.A(G57gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G85gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n320_), .B(new_n333_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n312_), .A2(KEYINPUT29), .ZN(new_n336_));
  XOR2_X1   g135(.A(G22gat), .B(G50gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT28), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n336_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n336_), .A2(new_n338_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n338_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(KEYINPUT92), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n262_), .B1(new_n312_), .B2(KEYINPUT29), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT91), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n218_), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n346_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n352_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n345_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n350_), .A2(new_n352_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n350_), .A2(new_n352_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n356_), .A2(new_n357_), .A3(new_n344_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT30), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n265_), .A2(KEYINPUT30), .A3(new_n266_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G227gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT85), .ZN(new_n367_));
  XOR2_X1   g166(.A(G71gat), .B(G99gat), .Z(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n362_), .A2(new_n363_), .A3(new_n360_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n365_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n369_), .B1(new_n373_), .B2(new_n364_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n315_), .B(KEYINPUT31), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT87), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n374_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n375_), .B(new_n376_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n359_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n344_), .B(new_n341_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n353_), .A2(new_n354_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n344_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n382_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n379_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n335_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n287_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT99), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n264_), .A2(new_n273_), .ZN(new_n393_));
  OAI221_X1 g192(.A(new_n335_), .B1(new_n283_), .B2(new_n392_), .C1(new_n393_), .C2(new_n391_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n334_), .A2(new_n395_), .ZN(new_n396_));
  OAI221_X1 g195(.A(new_n331_), .B1(new_n317_), .B2(new_n324_), .C1(new_n322_), .C2(new_n319_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n334_), .A2(new_n395_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n398_), .A2(new_n284_), .A3(new_n281_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n380_), .A2(new_n382_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(new_n359_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n390_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT65), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT64), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT64), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT6), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G99gat), .A2(G106gat), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n406_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n411_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n409_), .A2(KEYINPUT6), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n407_), .A2(KEYINPUT64), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n408_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT65), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G85gat), .B(G92gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT8), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT8), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT66), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT9), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G85gat), .A3(G92gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n426_), .B2(new_n435_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT10), .B(G99gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(G106gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n420_), .A3(new_n414_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n433_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n425_), .A2(new_n427_), .B1(new_n431_), .B2(KEYINPUT8), .ZN(new_n443_));
  INV_X1    g242(.A(new_n441_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT66), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G71gat), .B(G78gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(G57gat), .B(G64gat), .Z(new_n447_));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G64gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n446_), .A3(KEYINPUT11), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n442_), .A2(new_n445_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n442_), .A2(new_n445_), .A3(KEYINPUT67), .A4(new_n456_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n433_), .A2(new_n441_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n454_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT12), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(G230gat), .A2(G233gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n443_), .A2(new_n444_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(new_n454_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n459_), .A2(new_n460_), .A3(new_n464_), .A4(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n461_), .A2(new_n462_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n466_), .A2(new_n454_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n465_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G120gat), .B(G148gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G204gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT5), .B(G176gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  AND3_X1   g274(.A1(new_n468_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT68), .ZN(new_n478_));
  OAI22_X1  g277(.A1(new_n476_), .A2(new_n477_), .B1(new_n478_), .B2(KEYINPUT13), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n468_), .A2(new_n471_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n475_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n468_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n479_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G36gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G29gat), .ZN(new_n488_));
  INV_X1    g287(.A(G29gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G36gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G50gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G43gat), .ZN(new_n493_));
  INV_X1    g292(.A(G43gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G50gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n488_), .A2(new_n490_), .A3(new_n493_), .A4(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT15), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G1gat), .A2(G8gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT14), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G15gat), .A2(G22gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(G15gat), .A2(G22gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(G1gat), .ZN(new_n506_));
  INV_X1    g305(.A(G8gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n501_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n511_), .A2(new_n501_), .A3(new_n508_), .A4(new_n502_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n500_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n498_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n488_), .A2(new_n490_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n510_), .B(new_n512_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n499_), .A2(KEYINPUT77), .A3(new_n510_), .A4(new_n512_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n514_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT80), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT79), .ZN(new_n526_));
  INV_X1    g325(.A(new_n499_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n513_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n521_), .A2(KEYINPUT78), .A3(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n522_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n526_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  AOI221_X4 g334(.A(new_n530_), .B1(new_n527_), .B2(new_n513_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT78), .B1(new_n521_), .B2(new_n528_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n526_), .B(new_n534_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n525_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(G169gat), .ZN(new_n542_));
  INV_X1    g341(.A(G197gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n525_), .B(new_n544_), .C1(new_n535_), .C2(new_n539_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n486_), .A2(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n405_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n442_), .A2(new_n445_), .A3(new_n500_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n466_), .A2(new_n499_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT70), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT72), .A4(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT36), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(new_n557_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n551_), .A2(new_n552_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n558_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n551_), .B2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n559_), .B(new_n563_), .C1(new_n565_), .C2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT73), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n551_), .A2(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n558_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n551_), .A2(new_n552_), .A3(new_n564_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT73), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n559_), .A4(new_n563_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n559_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n570_), .A2(new_n576_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT37), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT75), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(new_n585_), .A3(new_n569_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n569_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n583_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n452_), .A2(new_n513_), .A3(new_n453_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n513_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n594_));
  INV_X1    g393(.A(G231gat), .ZN(new_n595_));
  INV_X1    g394(.A(G233gat), .ZN(new_n596_));
  OAI22_X1  g395(.A1(new_n593_), .A2(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n594_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n595_), .A2(new_n596_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(new_n592_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT16), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G183gat), .ZN(new_n605_));
  INV_X1    g404(.A(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n597_), .A2(new_n600_), .A3(KEYINPUT76), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n605_), .B(G211gat), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n601_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n608_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n591_), .A2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n550_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n506_), .A3(new_n335_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n588_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n614_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n550_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n335_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n620_), .A2(new_n621_), .A3(new_n627_), .ZN(G1324gat));
  INV_X1    g427(.A(new_n287_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n617_), .A2(new_n507_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  INV_X1    g430(.A(new_n625_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n629_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n633_), .B2(G8gat), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT39), .B(new_n507_), .C1(new_n632_), .C2(new_n629_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(new_n402_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G15gat), .B1(new_n625_), .B2(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT102), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT102), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(KEYINPUT41), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT41), .B1(new_n641_), .B2(new_n642_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n617_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(G15gat), .A3(new_n639_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n646_), .ZN(G1326gat));
  OAI21_X1  g446(.A(G22gat), .B1(new_n625_), .B2(new_n386_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n386_), .A2(G22gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n645_), .B2(new_n650_), .ZN(G1327gat));
  NAND2_X1  g450(.A1(new_n549_), .A2(new_n615_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n405_), .A2(new_n653_), .A3(new_n591_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n287_), .A2(new_n389_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n583_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT43), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n652_), .B1(new_n654_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT44), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n658_), .A2(KEYINPUT44), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n626_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n655_), .A2(new_n622_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n652_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n335_), .A2(new_n489_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT103), .Z(new_n667_));
  OAI22_X1  g466(.A1(new_n662_), .A2(new_n489_), .B1(new_n665_), .B2(new_n667_), .ZN(G1328gat));
  NOR2_X1   g467(.A1(new_n661_), .A2(new_n287_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n487_), .B1(new_n669_), .B2(new_n659_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n663_), .A2(new_n487_), .A3(new_n629_), .A4(new_n664_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT45), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n672_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n670_), .A2(new_n671_), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n671_), .B1(new_n670_), .B2(new_n676_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  INV_X1    g478(.A(KEYINPUT47), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n494_), .B1(new_n665_), .B2(new_n639_), .ZN(new_n682_));
  OAI211_X1 g481(.A(G43gat), .B(new_n402_), .C1(new_n658_), .C2(KEYINPUT44), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n681_), .B(new_n682_), .C1(new_n660_), .C2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n654_), .A2(new_n657_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n664_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n689_), .A2(G43gat), .A3(new_n402_), .A4(new_n659_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n681_), .B1(new_n690_), .B2(new_n682_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n680_), .B1(new_n685_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n682_), .B1(new_n660_), .B2(new_n683_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT106), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(KEYINPUT47), .A3(new_n684_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1330gat));
  NOR3_X1   g495(.A1(new_n661_), .A2(new_n492_), .A3(new_n386_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n663_), .A2(new_n359_), .A3(new_n664_), .ZN(new_n698_));
  AOI22_X1  g497(.A1(new_n697_), .A2(new_n659_), .B1(new_n492_), .B2(new_n698_), .ZN(G1331gat));
  NOR3_X1   g498(.A1(new_n655_), .A2(new_n548_), .A3(new_n486_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n624_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n626_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n616_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n335_), .A2(new_n328_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(G1332gat));
  OAI21_X1  g504(.A(G64gat), .B1(new_n701_), .B2(new_n287_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n287_), .A2(G64gat), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT108), .Z(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n703_), .B2(new_n710_), .ZN(G1333gat));
  OAI21_X1  g510(.A(G71gat), .B1(new_n701_), .B2(new_n639_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT49), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n639_), .A2(G71gat), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT109), .Z(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n703_), .B2(new_n715_), .ZN(G1334gat));
  OAI21_X1  g515(.A(G78gat), .B1(new_n701_), .B2(new_n386_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT50), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n386_), .A2(G78gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n703_), .B2(new_n719_), .ZN(G1335gat));
  NOR2_X1   g519(.A1(new_n486_), .A2(new_n548_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n615_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n654_), .B2(new_n657_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n626_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n663_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1336gat));
  OAI21_X1  g529(.A(G92gat), .B1(new_n724_), .B2(new_n287_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n205_), .A3(new_n629_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1337gat));
  INV_X1    g532(.A(G99gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n723_), .B2(new_n402_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n727_), .A2(new_n438_), .A3(new_n639_), .ZN(new_n736_));
  OAI22_X1  g535(.A1(new_n735_), .A2(new_n736_), .B1(KEYINPUT110), .B2(KEYINPUT51), .ZN(new_n737_));
  NAND2_X1  g536(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT111), .Z(new_n739_));
  XNOR2_X1  g538(.A(new_n737_), .B(new_n739_), .ZN(G1338gat));
  INV_X1    g539(.A(G106gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n723_), .B2(new_n359_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT52), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(KEYINPUT52), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n663_), .A2(new_n741_), .A3(new_n359_), .A4(new_n726_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT112), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g547(.A1(new_n548_), .A2(G113gat), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT120), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT59), .ZN(new_n751_));
  INV_X1    g550(.A(new_n469_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n459_), .A2(new_n752_), .A3(new_n460_), .A4(new_n464_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n465_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n468_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n463_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n757_), .A2(KEYINPUT55), .A3(new_n460_), .A4(new_n467_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n481_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT56), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n481_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n533_), .A2(new_n522_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n514_), .A2(new_n521_), .A3(new_n534_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n545_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n547_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(new_n476_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(KEYINPUT58), .A3(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n481_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n481_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n591_), .A2(new_n770_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n476_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n768_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n586_), .A2(KEYINPUT57), .A3(new_n587_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT118), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n785_), .B(new_n782_), .C1(new_n778_), .C2(new_n780_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n776_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n588_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n789_));
  XOR2_X1   g588(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n790_));
  OAI21_X1  g589(.A(new_n788_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n790_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n779_), .B1(new_n764_), .B2(new_n777_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT117), .B(new_n792_), .C1(new_n793_), .C2(new_n588_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n615_), .B1(new_n787_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n546_), .A2(new_n614_), .A3(new_n547_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n546_), .A2(new_n614_), .A3(KEYINPUT113), .A4(new_n547_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n797_), .B1(new_n802_), .B2(new_n486_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n486_), .A2(new_n797_), .A3(new_n800_), .A4(new_n801_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n656_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT115), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n479_), .A2(new_n485_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n800_), .A2(new_n801_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT114), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n804_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n656_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n807_), .A2(KEYINPUT54), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n811_), .A2(new_n812_), .A3(new_n656_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n812_), .B1(new_n811_), .B2(new_n656_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n796_), .A2(new_n814_), .A3(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n402_), .A2(new_n335_), .A3(new_n386_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n629_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n751_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n751_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n816_), .A2(new_n817_), .A3(new_n815_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT54), .B1(new_n807_), .B2(new_n813_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n789_), .A2(new_n790_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n615_), .B1(new_n787_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n823_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n750_), .B1(new_n822_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n828_), .A2(new_n814_), .A3(new_n818_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n751_), .A3(new_n821_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n821_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n826_), .B2(new_n796_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT120), .B(new_n832_), .C1(new_n834_), .C2(new_n751_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n749_), .B1(new_n830_), .B2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n819_), .A2(new_n548_), .A3(new_n821_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n837_), .A2(KEYINPUT119), .A3(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n836_), .A2(new_n843_), .ZN(G1340gat));
  NOR3_X1   g643(.A1(new_n822_), .A2(new_n829_), .A3(new_n486_), .ZN(new_n845_));
  INV_X1    g644(.A(G120gat), .ZN(new_n846_));
  INV_X1    g645(.A(new_n834_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n486_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(KEYINPUT60), .B2(new_n846_), .ZN(new_n849_));
  OAI22_X1  g648(.A1(new_n845_), .A2(new_n846_), .B1(new_n847_), .B2(new_n849_), .ZN(G1341gat));
  AOI21_X1  g649(.A(G127gat), .B1(new_n834_), .B2(new_n614_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n830_), .A2(new_n835_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n614_), .A2(G127gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1342gat));
  AOI21_X1  g653(.A(G134gat), .B1(new_n834_), .B2(new_n588_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n591_), .A2(G134gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n852_), .B2(new_n856_), .ZN(G1343gat));
  INV_X1    g656(.A(new_n819_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n629_), .A2(new_n626_), .A3(new_n383_), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(KEYINPUT121), .Z(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n548_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n808_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT122), .B(G148gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1345gat));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n614_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT123), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n867_), .B(new_n869_), .ZN(G1346gat));
  INV_X1    g669(.A(G162gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n861_), .A2(new_n871_), .A3(new_n588_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n861_), .A2(new_n591_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n874_), .B2(new_n871_), .ZN(G1347gat));
  NAND2_X1  g674(.A1(new_n629_), .A2(new_n626_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n639_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n359_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n831_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n548_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G169gat), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n880_), .A2(new_n548_), .A3(new_n241_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n881_), .A2(G169gat), .A3(new_n883_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .ZN(G1348gat));
  NAND2_X1  g687(.A1(new_n880_), .A2(new_n808_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n858_), .A2(new_n359_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n878_), .A2(new_n222_), .A3(new_n486_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n889_), .A2(new_n238_), .B1(new_n890_), .B2(new_n891_), .ZN(G1349gat));
  INV_X1    g691(.A(new_n880_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n893_), .A2(new_n251_), .A3(new_n615_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(new_n614_), .A3(new_n877_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n229_), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n893_), .B2(new_n656_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n880_), .A2(new_n228_), .A3(new_n588_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1351gat));
  NOR2_X1   g698(.A1(new_n876_), .A2(new_n383_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n819_), .A2(new_n548_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n543_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n901_), .B2(new_n543_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n901_), .A2(new_n543_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(G1352gat));
  AND2_X1   g705(.A1(new_n819_), .A2(new_n900_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n808_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g708(.A(new_n615_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT126), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n911_), .B(new_n913_), .ZN(G1354gat));
  NAND2_X1  g713(.A1(new_n907_), .A2(new_n588_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT127), .B(G218gat), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n656_), .A2(new_n916_), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n915_), .A2(new_n916_), .B1(new_n907_), .B2(new_n917_), .ZN(G1355gat));
endmodule


