//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G120gat), .B(G148gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT5), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G176gat), .B(G204gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  XNOR2_X1  g006(.A(G57gat), .B(G64gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n210_));
  XOR2_X1   g009(.A(G71gat), .B(G78gat), .Z(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n210_), .A2(new_n211_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G85gat), .B(G92gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT7), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n217_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT8), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(new_n217_), .C1(new_n220_), .C2(new_n223_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n221_), .B(KEYINPUT6), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT9), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT66), .B(G85gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(G92gat), .ZN(new_n232_));
  OAI221_X1 g031(.A(new_n229_), .B1(new_n230_), .B2(new_n216_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n236_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n234_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT10), .B(G99gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT64), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT65), .A3(new_n234_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n233_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n228_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n231_), .A2(new_n232_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n216_), .A2(new_n230_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n251_), .A2(new_n252_), .A3(new_n223_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT65), .B1(new_n246_), .B2(new_n234_), .ZN(new_n254_));
  AOI211_X1 g053(.A(new_n241_), .B(G106gat), .C1(new_n244_), .C2(new_n245_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(KEYINPUT67), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n215_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(KEYINPUT67), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n248_), .A2(new_n249_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(new_n228_), .A4(new_n214_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n258_), .A2(KEYINPUT12), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n263_), .B(new_n215_), .C1(new_n250_), .C2(new_n257_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT68), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n266_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n268_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n203_), .B(new_n207_), .C1(new_n270_), .C2(new_n274_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n272_), .A2(new_n207_), .A3(new_n268_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n207_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n267_), .A2(KEYINPUT68), .A3(new_n269_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n273_), .B1(new_n272_), .B2(new_n268_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(new_n203_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n202_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n276_), .B1(new_n282_), .B2(new_n203_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n207_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT69), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(KEYINPUT13), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291_));
  INV_X1    g090(.A(G1gat), .ZN(new_n292_));
  INV_X1    g091(.A(G8gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT14), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G8gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n214_), .B(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G127gat), .B(G155gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT16), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G183gat), .B(G211gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT17), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n304_), .A2(new_n305_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n300_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(new_n306_), .B2(new_n300_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT76), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G190gat), .B(G218gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT72), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G134gat), .B(G162gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT36), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G29gat), .B(G36gat), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT70), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(KEYINPUT70), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G43gat), .B(G50gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT15), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(KEYINPUT15), .A3(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n330_));
  INV_X1    g129(.A(new_n324_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n259_), .A2(new_n260_), .A3(new_n331_), .A4(new_n228_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G232gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT34), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT35), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .A4(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n336_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n329_), .A2(new_n332_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n337_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n329_), .B2(KEYINPUT71), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n338_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n315_), .B1(new_n343_), .B2(KEYINPUT74), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n345_), .B(new_n338_), .C1(new_n340_), .C2(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n314_), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n343_), .B2(new_n315_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT37), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n310_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n290_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT77), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  INV_X1    g157(.A(G43gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(G15gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n360_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366_));
  INV_X1    g165(.A(G169gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(KEYINPUT22), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369_));
  AOI21_X1  g168(.A(G176gat), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT22), .B1(new_n367_), .B2(KEYINPUT80), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n366_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT22), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n373_), .A3(G169gat), .ZN(new_n374_));
  INV_X1    g173(.A(G176gat), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n371_), .A2(new_n374_), .A3(new_n366_), .A4(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n365_), .B1(new_n372_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT23), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT79), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT23), .ZN(new_n383_));
  AND2_X1   g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n387_), .B2(KEYINPUT23), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .A4(new_n386_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT84), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n371_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT81), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n396_), .A2(KEYINPUT82), .A3(new_n377_), .A4(new_n376_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n389_), .A2(new_n398_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n379_), .A2(new_n394_), .A3(new_n397_), .A4(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n387_), .A2(KEYINPUT23), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n381_), .A2(new_n383_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(new_n387_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT25), .B(G183gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT26), .B(G190gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT78), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(G169gat), .B2(G176gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT24), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n410_), .A3(new_n377_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n406_), .B(new_n413_), .C1(new_n412_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n400_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n364_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G127gat), .B(G134gat), .Z(new_n421_));
  XOR2_X1   g220(.A(G113gat), .B(G120gat), .Z(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT31), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n418_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n416_), .B(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT85), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n420_), .B(new_n424_), .C1(new_n429_), .C2(new_n363_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n424_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n363_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n419_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G155gat), .A2(G162gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n439_));
  NOR4_X1   g238(.A1(new_n439_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT87), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G141gat), .A2(G148gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT2), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT2), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G141gat), .A3(G148gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(G141gat), .A2(G148gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT3), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n444_), .A2(new_n452_), .A3(KEYINPUT88), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n439_), .B1(new_n450_), .B2(KEYINPUT3), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n441_), .A2(KEYINPUT87), .A3(new_n442_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n446_), .A2(new_n448_), .B1(new_n450_), .B2(KEYINPUT3), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n454_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n438_), .B1(new_n453_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n423_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n437_), .B1(KEYINPUT1), .B2(new_n435_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(KEYINPUT1), .B2(new_n435_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n450_), .A3(new_n445_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n438_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT88), .B1(new_n444_), .B2(new_n452_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(new_n458_), .A3(new_n454_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n464_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n423_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n465_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n465_), .A2(new_n471_), .A3(KEYINPUT4), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n475_), .B(new_n423_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n472_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n473_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G29gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G57gat), .B(G85gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n479_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n473_), .B(new_n484_), .C1(new_n474_), .C2(new_n478_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G22gat), .B(G50gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n469_), .A2(new_n470_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n490_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n490_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502_));
  INV_X1    g301(.A(G218gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G211gat), .ZN(new_n504_));
  INV_X1    g303(.A(G211gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G218gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n502_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G197gat), .B(G204gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT21), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n504_), .A2(new_n506_), .A3(new_n502_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n508_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n510_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n512_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n507_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n517_));
  INV_X1    g316(.A(G204gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(G197gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT21), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(KEYINPUT91), .B2(new_n509_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n513_), .B1(new_n516_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(KEYINPUT90), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G228gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT89), .ZN(new_n527_));
  INV_X1    g326(.A(G78gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n234_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n530_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n501_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n497_), .A2(new_n500_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G226gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT19), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n523_), .B1(new_n400_), .B2(new_n415_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n377_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT22), .B(G169gat), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n541_), .B2(new_n375_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n403_), .B2(new_n390_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n404_), .A2(new_n405_), .ZN(new_n544_));
  AND2_X1   g343(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n545_));
  NOR2_X1   g344(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n407_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n389_), .A2(new_n544_), .A3(new_n548_), .A4(new_n392_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n414_), .A2(new_n547_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n543_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT20), .B1(new_n551_), .B2(new_n522_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n538_), .B1(new_n539_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n400_), .A2(new_n523_), .A3(new_n415_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n538_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n551_), .B2(new_n522_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G64gat), .B(G92gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(G8gat), .A2(G36gat), .ZN(new_n562_));
  NOR2_X1   g361(.A1(G8gat), .A2(G36gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n566_));
  INV_X1    g365(.A(G92gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G64gat), .ZN(new_n568_));
  INV_X1    g367(.A(G64gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(G92gat), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n568_), .B(new_n570_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n565_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n566_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G8gat), .B(G36gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(new_n560_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n571_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n573_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n559_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n554_), .A2(new_n557_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n538_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n416_), .A2(new_n522_), .ZN(new_n581_));
  OAI211_X1 g380(.A(KEYINPUT20), .B(new_n555_), .C1(new_n551_), .C2(new_n522_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n572_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n580_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n578_), .A2(KEYINPUT27), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n580_), .A2(new_n584_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT27), .B1(new_n589_), .B2(new_n586_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n434_), .A2(new_n489_), .A3(new_n536_), .A4(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n534_), .A2(new_n535_), .A3(new_n487_), .A4(new_n486_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n593_), .A2(new_n587_), .A3(new_n590_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n487_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n465_), .A2(new_n471_), .A3(KEYINPUT4), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n477_), .A3(new_n476_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n484_), .B1(new_n597_), .B2(new_n473_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n585_), .B2(KEYINPUT32), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT32), .ZN(new_n601_));
  AOI211_X1 g400(.A(KEYINPUT96), .B(new_n601_), .C1(new_n577_), .C2(new_n572_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT97), .B1(new_n604_), .B2(new_n580_), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n539_), .A2(new_n582_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n555_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  OAI22_X1  g408(.A1(new_n595_), .A2(new_n598_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n585_), .A2(KEYINPUT32), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT98), .B1(new_n559_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n614_), .B(new_n611_), .C1(new_n553_), .C2(new_n558_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT99), .B1(new_n610_), .B2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n611_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT98), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n604_), .A2(KEYINPUT97), .A3(new_n580_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n608_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n486_), .A2(new_n487_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n595_), .A2(KEYINPUT33), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n596_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n465_), .A2(new_n471_), .A3(new_n477_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(new_n485_), .ZN(new_n629_));
  AOI22_X1  g428(.A1(new_n487_), .A2(new_n626_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n625_), .A2(new_n630_), .A3(new_n586_), .A4(new_n589_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n617_), .A2(new_n624_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n594_), .B1(new_n632_), .B2(new_n536_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT86), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n434_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n430_), .A2(new_n433_), .A3(KEYINPUT86), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n592_), .B1(new_n633_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n328_), .A2(new_n297_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n324_), .A2(new_n297_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n324_), .B(new_n297_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G113gat), .B(G141gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G169gat), .B(G197gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(new_n649_));
  XNOR2_X1  g448(.A(new_n646_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n638_), .A2(KEYINPUT100), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n638_), .B2(new_n651_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n357_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n488_), .A2(new_n292_), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n284_), .A2(new_n288_), .A3(new_n651_), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n658_), .A2(KEYINPUT101), .A3(new_n310_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT101), .B1(new_n658_), .B2(new_n310_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n347_), .A2(new_n350_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n638_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n489_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n655_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n657_), .A2(new_n664_), .A3(new_n665_), .ZN(G1324gat));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  INV_X1    g466(.A(new_n663_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n591_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n667_), .B1(new_n670_), .B2(G8gat), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT39), .B(new_n293_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n293_), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n671_), .A2(new_n672_), .B1(new_n654_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g474(.A(new_n637_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G15gat), .B1(new_n663_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n678_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n676_), .A2(G15gat), .ZN(new_n681_));
  OAI22_X1  g480(.A1(new_n679_), .A2(new_n680_), .B1(new_n654_), .B2(new_n681_), .ZN(G1326gat));
  XNOR2_X1  g481(.A(new_n536_), .B(KEYINPUT102), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G22gat), .B1(new_n663_), .B2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n684_), .A2(G22gat), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n686_), .A2(new_n687_), .B1(new_n654_), .B2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n310_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n289_), .A2(new_n690_), .A3(new_n661_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n691_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT104), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n694_), .B(new_n691_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(G29gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n488_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n658_), .A2(KEYINPUT103), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n352_), .A2(new_n354_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n638_), .A2(KEYINPUT43), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT43), .B1(new_n638_), .B2(new_n702_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n690_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n699_), .B(new_n700_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n638_), .A2(new_n702_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n638_), .A2(KEYINPUT43), .A3(new_n702_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n310_), .A3(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(KEYINPUT103), .B(KEYINPUT44), .C1(new_n712_), .C2(new_n658_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n489_), .B1(new_n707_), .B2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n698_), .B1(new_n714_), .B2(new_n697_), .ZN(G1328gat));
  NOR2_X1   g514(.A1(new_n591_), .A2(G36gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n693_), .A2(new_n695_), .A3(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT106), .B(KEYINPUT108), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n717_), .B(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n707_), .A2(new_n713_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(KEYINPUT105), .A3(new_n669_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT105), .B1(new_n722_), .B2(new_n669_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT46), .B(new_n721_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  NAND2_X1  g529(.A1(new_n696_), .A2(new_n637_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n359_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n434_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n359_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n722_), .A2(KEYINPUT109), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT109), .B1(new_n722_), .B2(new_n734_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT47), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n732_), .B(new_n739_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n696_), .B2(new_n683_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n536_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(G50gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n722_), .B2(new_n744_), .ZN(G1331gat));
  NOR2_X1   g544(.A1(new_n290_), .A2(new_n651_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n690_), .A3(new_n662_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G57gat), .B1(new_n747_), .B2(new_n489_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n746_), .A2(new_n638_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(new_n355_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n489_), .A2(G57gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT110), .ZN(G1332gat));
  NAND3_X1  g553(.A1(new_n750_), .A2(new_n569_), .A3(new_n669_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G64gat), .B1(new_n747_), .B2(new_n591_), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n757_));
  OR2_X1    g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n756_), .A2(new_n757_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n759_), .B2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n747_), .B2(new_n676_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n676_), .A2(G71gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n751_), .B2(new_n764_), .ZN(G1334gat));
  NAND3_X1  g564(.A1(new_n750_), .A2(new_n528_), .A3(new_n683_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G78gat), .B1(new_n747_), .B2(new_n684_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n767_), .A2(new_n768_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n766_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  NAND2_X1  g571(.A1(new_n705_), .A2(new_n746_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n773_), .A2(new_n489_), .A3(new_n231_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n661_), .ZN(new_n775_));
  AND4_X1   g574(.A1(new_n638_), .A2(new_n746_), .A3(new_n310_), .A4(new_n775_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(new_n488_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n777_), .A2(G85gat), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n778_), .A2(KEYINPUT113), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(KEYINPUT113), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n774_), .B1(new_n779_), .B2(new_n780_), .ZN(G1336gat));
  OAI21_X1  g580(.A(G92gat), .B1(new_n773_), .B2(new_n591_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n567_), .A3(new_n669_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1337gat));
  NAND3_X1  g583(.A1(new_n776_), .A2(new_n434_), .A3(new_n246_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT114), .ZN(new_n786_));
  OAI21_X1  g585(.A(G99gat), .B1(new_n773_), .B2(new_n676_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n776_), .A2(new_n234_), .A3(new_n743_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n746_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n712_), .A2(new_n536_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n234_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT115), .B1(new_n773_), .B2(new_n536_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n790_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n790_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  NAND4_X1  g602(.A1(new_n284_), .A2(new_n288_), .A3(new_n355_), .A4(new_n650_), .ZN(new_n804_));
  XOR2_X1   g603(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n651_), .A2(new_n277_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n262_), .A2(new_n271_), .A3(new_n264_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT55), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n267_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n265_), .A2(KEYINPUT55), .A3(new_n266_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n272_), .A2(KEYINPUT117), .A3(KEYINPUT55), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n207_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n207_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n809_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n639_), .A2(new_n640_), .A3(new_n644_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n649_), .B1(new_n643_), .B2(new_n641_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n825_), .A2(KEYINPUT118), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(KEYINPUT118), .ZN(new_n827_));
  INV_X1    g626(.A(new_n649_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n826_), .B(new_n827_), .C1(new_n646_), .C2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n661_), .B1(new_n822_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n829_), .A2(new_n276_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n207_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n207_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n701_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT58), .B(new_n834_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT57), .B(new_n661_), .C1(new_n822_), .C2(new_n830_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n833_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n808_), .B1(new_n843_), .B2(new_n310_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n743_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n733_), .A2(new_n489_), .A3(new_n669_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n651_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n651_), .A2(G113gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT119), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n849_), .B1(new_n853_), .B2(new_n855_), .ZN(G1340gat));
  XNOR2_X1  g655(.A(KEYINPUT120), .B(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n290_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n848_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n857_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n290_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n857_), .ZN(G1341gat));
  INV_X1    g660(.A(G127gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n848_), .A2(new_n862_), .A3(new_n690_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n310_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n848_), .A2(new_n866_), .A3(new_n775_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n701_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n866_), .ZN(G1343gat));
  NOR4_X1   g668(.A1(new_n637_), .A2(new_n489_), .A3(new_n536_), .A4(new_n669_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT121), .B1(new_n844_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n832_), .A2(new_n831_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n690_), .B1(new_n874_), .B2(new_n842_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n873_), .B(new_n870_), .C1(new_n875_), .C2(new_n808_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n651_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n289_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n690_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT61), .B(G155gat), .Z(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n885_));
  INV_X1    g684(.A(new_n883_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n877_), .A2(new_n690_), .A3(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(new_n885_), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n885_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n886_), .B1(new_n877_), .B2(new_n690_), .ZN(new_n890_));
  AOI211_X1 g689(.A(new_n310_), .B(new_n883_), .C1(new_n872_), .C2(new_n876_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1346gat));
  INV_X1    g692(.A(new_n877_), .ZN(new_n894_));
  OR3_X1    g693(.A1(new_n894_), .A2(G162gat), .A3(new_n661_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G162gat), .B1(new_n894_), .B2(new_n701_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1347gat));
  NOR3_X1   g696(.A1(new_n676_), .A2(new_n488_), .A3(new_n591_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n684_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n844_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n367_), .B1(new_n900_), .B2(new_n651_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n901_), .A2(KEYINPUT62), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n541_), .A3(new_n651_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(KEYINPUT62), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(G1348gat));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n844_), .B2(new_n743_), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT124), .B(new_n536_), .C1(new_n875_), .C2(new_n808_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n898_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n909_), .A2(new_n375_), .A3(new_n290_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G176gat), .B1(new_n900_), .B2(new_n289_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1349gat));
  INV_X1    g711(.A(G183gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n909_), .B2(new_n310_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n900_), .ZN(new_n915_));
  OR3_X1    g714(.A1(new_n915_), .A2(new_n404_), .A3(new_n310_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n914_), .A2(new_n916_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n915_), .B2(new_n701_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n900_), .A2(new_n405_), .A3(new_n775_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1351gat));
  NOR4_X1   g723(.A1(new_n844_), .A2(new_n593_), .A3(new_n591_), .A4(new_n637_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n651_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n289_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT126), .B(G204gat), .Z(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1353gat));
  AOI21_X1  g729(.A(new_n310_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n925_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT127), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n925_), .A2(new_n934_), .A3(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n933_), .A2(new_n935_), .A3(new_n937_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1354gat));
  NAND3_X1  g740(.A1(new_n925_), .A2(new_n503_), .A3(new_n775_), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n925_), .A2(new_n702_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n503_), .ZN(G1355gat));
endmodule


