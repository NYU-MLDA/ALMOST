//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  NAND3_X1  g001(.A1(new_n202_), .A2(G183gat), .A3(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND4_X1  g004(.A1(new_n202_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT83), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT23), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n207_), .B2(KEYINPUT23), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n205_), .B(new_n206_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n212_), .A2(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n215_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n222_));
  AOI21_X1  g021(.A(G176gat), .B1(new_n222_), .B2(KEYINPUT85), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT86), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT22), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT86), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n227_), .A3(G169gat), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n226_), .A2(KEYINPUT85), .A3(G169gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n203_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n218_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n220_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G15gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT31), .Z(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n245_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n241_), .B(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(G233gat), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT94), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  AND2_X1   g055(.A1(G197gat), .A2(G204gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G197gat), .A2(G204gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n256_), .A2(KEYINPUT95), .ZN(new_n260_));
  OR2_X1    g059(.A1(G197gat), .A2(G204gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G197gat), .A2(G204gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G218gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G211gat), .ZN(new_n265_));
  INV_X1    g064(.A(G211gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G218gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n259_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G211gat), .B(G218gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n257_), .A2(new_n258_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n260_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT88), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G155gat), .A3(G162gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT89), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n275_), .A2(new_n277_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT1), .ZN(new_n289_));
  INV_X1    g088(.A(new_n282_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n279_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT89), .ZN(new_n292_));
  INV_X1    g091(.A(new_n286_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT90), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n297_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n285_), .A2(new_n300_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n302_));
  AND3_X1   g101(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n299_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n282_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT91), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT91), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n287_), .A2(new_n294_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n255_), .B(new_n273_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n282_), .B1(new_n288_), .B2(KEYINPUT1), .ZN(new_n314_));
  AOI211_X1 g113(.A(KEYINPUT89), .B(new_n286_), .C1(new_n314_), .C2(new_n279_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n292_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n305_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n309_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n318_));
  OAI22_X1  g117(.A1(new_n315_), .A2(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT96), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n263_), .A2(new_n268_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n271_), .A2(new_n270_), .A3(new_n260_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(KEYINPUT96), .A4(new_n259_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n319_), .A2(KEYINPUT29), .B1(new_n321_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n313_), .B1(new_n255_), .B2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n311_), .A2(new_n312_), .A3(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n319_), .B2(KEYINPUT29), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G78gat), .B(G106gat), .Z(new_n332_));
  XNOR2_X1  g131(.A(G22gat), .B(G50gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n330_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n335_), .B(new_n313_), .C1(new_n255_), .C2(new_n325_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n331_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n319_), .A2(KEYINPUT100), .A3(new_n248_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n287_), .A2(new_n294_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n308_), .A2(new_n310_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n248_), .A2(KEYINPUT100), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n248_), .A2(KEYINPUT100), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .A4(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT101), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n248_), .A2(KEYINPUT4), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n348_), .B1(new_n311_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n350_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n346_), .A2(KEYINPUT4), .ZN(new_n360_));
  INV_X1    g159(.A(new_n354_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n355_), .A2(new_n359_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365_));
  XOR2_X1   g164(.A(G8gat), .B(G36gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n321_), .A2(new_n220_), .A3(new_n236_), .A4(new_n324_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n226_), .A2(G169gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n222_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n218_), .B1(new_n374_), .B2(G176gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n211_), .B2(new_n234_), .ZN(new_n376_));
  INV_X1    g175(.A(G183gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT25), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G183gat), .ZN(new_n380_));
  INV_X1    g179(.A(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT26), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT26), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G190gat), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n378_), .A2(new_n380_), .A3(new_n382_), .A4(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n215_), .A2(new_n214_), .ZN(new_n386_));
  AND4_X1   g185(.A1(new_n219_), .A2(new_n385_), .A3(new_n386_), .A4(new_n232_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n273_), .B1(new_n376_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n372_), .A2(new_n388_), .A3(KEYINPUT20), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n390_));
  AND2_X1   g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n322_), .A2(new_n323_), .A3(new_n259_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n216_), .A2(new_n219_), .A3(new_n232_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n205_), .A2(new_n206_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n210_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT23), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n233_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n393_), .B(new_n394_), .C1(new_n399_), .C2(new_n375_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT98), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n376_), .A2(new_n387_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT98), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n393_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n321_), .A2(new_n324_), .ZN(new_n407_));
  AOI211_X1 g206(.A(new_n406_), .B(new_n392_), .C1(new_n407_), .C2(new_n237_), .ZN(new_n408_));
  AOI221_X4 g207(.A(new_n371_), .B1(new_n389_), .B2(new_n392_), .C1(new_n405_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n392_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT103), .B(new_n394_), .C1(new_n399_), .C2(new_n375_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT103), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n376_), .B2(new_n387_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(new_n393_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n406_), .B1(new_n407_), .B2(new_n237_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT104), .ZN(new_n417_));
  OAI22_X1  g216(.A1(new_n416_), .A2(new_n417_), .B1(new_n392_), .B2(new_n389_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n416_), .A2(new_n417_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n371_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n409_), .B1(new_n420_), .B2(KEYINPUT106), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT106), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n422_), .B(new_n371_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n365_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n403_), .B1(new_n402_), .B2(new_n393_), .ZN(new_n425_));
  NOR4_X1   g224(.A1(new_n376_), .A2(new_n273_), .A3(new_n387_), .A4(KEYINPUT98), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n410_), .B(new_n415_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n389_), .A2(new_n392_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n370_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n409_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n365_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n339_), .B(new_n364_), .C1(new_n424_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  INV_X1    g233(.A(new_n359_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n350_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n352_), .A2(new_n354_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n434_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT102), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n346_), .A2(new_n348_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n349_), .B1(new_n311_), .B2(new_n353_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n441_), .B(new_n359_), .C1(new_n352_), .C2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n430_), .A2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n350_), .B(new_n435_), .C1(new_n352_), .C2(new_n354_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT102), .A3(new_n434_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n362_), .A2(KEYINPUT33), .A3(new_n363_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n440_), .A2(new_n444_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n355_), .A2(new_n359_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n370_), .A2(KEYINPUT32), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n427_), .A2(new_n451_), .A3(new_n428_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n339_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n433_), .B1(new_n456_), .B2(KEYINPUT105), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT105), .ZN(new_n458_));
  AOI211_X1 g257(.A(new_n458_), .B(new_n339_), .C1(new_n448_), .C2(new_n455_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n250_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n424_), .A2(new_n432_), .ZN(new_n461_));
  NOR4_X1   g260(.A1(new_n461_), .A2(new_n250_), .A3(new_n339_), .A4(new_n450_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  INV_X1    g264(.A(G1gat), .ZN(new_n466_));
  INV_X1    g265(.A(G8gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n471_), .B(new_n474_), .Z(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(G229gat), .A3(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n474_), .B(KEYINPUT15), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n471_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n471_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n474_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT82), .Z(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G169gat), .B(G197gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n476_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n464_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G120gat), .B(G148gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT75), .ZN(new_n495_));
  XOR2_X1   g294(.A(G176gat), .B(G204gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT76), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n495_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  INV_X1    g299(.A(KEYINPUT73), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT77), .Z(new_n503_));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n504_));
  XOR2_X1   g303(.A(G85gat), .B(G92gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT66), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT8), .ZN(new_n508_));
  NOR2_X1   g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT7), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT6), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(G99gat), .A3(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n507_), .A2(new_n508_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT67), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n512_), .A2(new_n514_), .A3(KEYINPUT67), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n518_), .B1(new_n522_), .B2(KEYINPUT68), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT68), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n524_), .A3(new_n521_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n506_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n517_), .B1(new_n526_), .B2(new_n508_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n505_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT10), .B(G99gat), .Z(new_n529_));
  INV_X1    g328(.A(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT9), .ZN(new_n532_));
  INV_X1    g331(.A(G85gat), .ZN(new_n533_));
  INV_X1    g332(.A(G92gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n533_), .A2(new_n534_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT65), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n532_), .B(new_n535_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n528_), .A2(new_n531_), .A3(new_n515_), .A4(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n527_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT69), .B(G71gat), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n542_), .A2(G78gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(G78gat), .ZN(new_n544_));
  OAI211_X1 g343(.A(KEYINPUT11), .B(new_n541_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT69), .B(G71gat), .Z(new_n547_));
  INV_X1    g346(.A(G78gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n542_), .A2(G78gat), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n546_), .A2(new_n549_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n545_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n545_), .B2(new_n552_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n504_), .B1(new_n540_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n527_), .A2(new_n557_), .A3(new_n539_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT64), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n539_), .B(KEYINPUT72), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n527_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n556_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n504_), .B1(new_n566_), .B2(new_n554_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n558_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n559_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n557_), .B1(new_n527_), .B2(new_n539_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n561_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n503_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n502_), .B(KEYINPUT77), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(KEYINPUT13), .A3(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT79), .ZN(new_n585_));
  XOR2_X1   g384(.A(G134gat), .B(G162gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n540_), .A2(new_n474_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n565_), .A2(new_n477_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT34), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n592_), .B2(KEYINPUT78), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n590_), .B1(new_n594_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n593_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n589_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n594_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n593_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n589_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .A4(new_n590_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n604_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT37), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n557_), .B(new_n479_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT81), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT17), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n613_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT17), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n613_), .B1(new_n622_), .B2(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n583_), .A2(new_n610_), .A3(new_n624_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n493_), .A2(KEYINPUT107), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT107), .B1(new_n493_), .B2(new_n625_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n364_), .A2(G1gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT108), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT108), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n626_), .A2(new_n631_), .A3(new_n627_), .A4(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(KEYINPUT38), .A3(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n464_), .A2(new_n609_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n624_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n582_), .A2(new_n491_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n637_), .A2(new_n364_), .A3(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n635_), .B(new_n636_), .C1(new_n466_), .C2(new_n641_), .ZN(G1324gat));
  NAND4_X1  g441(.A1(new_n626_), .A2(new_n467_), .A3(new_n461_), .A4(new_n627_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n464_), .A2(new_n461_), .A3(new_n639_), .A4(new_n609_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT109), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n646_), .ZN(new_n649_));
  AND4_X1   g448(.A1(new_n644_), .A2(new_n648_), .A3(G8gat), .A4(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n647_), .A2(new_n467_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n644_), .B1(new_n651_), .B2(new_n649_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n643_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT40), .B(new_n643_), .C1(new_n650_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1325gat));
  INV_X1    g456(.A(G15gat), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n637_), .A2(new_n640_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n250_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT41), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n493_), .A2(new_n625_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n339_), .B(KEYINPUT110), .Z(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n659_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT42), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n663_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(new_n609_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n638_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n582_), .A2(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n464_), .A2(new_n492_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n450_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n582_), .A2(new_n491_), .A3(new_n624_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT37), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n609_), .B(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n464_), .B2(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT43), .B(new_n610_), .C1(new_n460_), .C2(new_n463_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT44), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n678_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n453_), .A2(new_n454_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n364_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n430_), .B(new_n443_), .C1(new_n445_), .C2(new_n434_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT102), .B1(new_n445_), .B2(new_n434_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n689_), .B1(new_n692_), .B2(new_n446_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n458_), .B1(new_n693_), .B2(new_n339_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n456_), .A2(KEYINPUT105), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n433_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n462_), .B1(new_n696_), .B2(new_n250_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n697_), .B2(new_n610_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n464_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n687_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT111), .ZN(new_n701_));
  AOI22_X1  g500(.A1(new_n686_), .A2(new_n701_), .B1(KEYINPUT44), .B2(new_n700_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n450_), .A2(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n677_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  AND2_X1   g503(.A1(new_n421_), .A2(new_n423_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n431_), .B1(new_n705_), .B2(new_n365_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(KEYINPUT112), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(KEYINPUT112), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n464_), .A2(new_n710_), .A3(new_n492_), .A4(new_n675_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(KEYINPUT113), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(KEYINPUT113), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n676_), .A2(new_n716_), .A3(new_n710_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n711_), .A2(KEYINPUT113), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT45), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n715_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT44), .B(new_n678_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n461_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n686_), .B2(new_n701_), .ZN(new_n723_));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT46), .B(new_n720_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n714_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n717_), .A2(new_n718_), .A3(KEYINPUT45), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(new_n700_), .B2(KEYINPUT111), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n685_), .B(new_n687_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n461_), .B(new_n721_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n728_), .B1(new_n732_), .B2(G36gat), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT114), .B(KEYINPUT46), .Z(new_n734_));
  OAI21_X1  g533(.A(new_n725_), .B1(new_n733_), .B2(new_n734_), .ZN(G1329gat));
  AND2_X1   g534(.A1(new_n660_), .A2(G43gat), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n721_), .B(new_n736_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT115), .B(G43gat), .Z(new_n738_));
  INV_X1    g537(.A(new_n676_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n250_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT47), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n737_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1330gat));
  INV_X1    g544(.A(new_n339_), .ZN(new_n746_));
  INV_X1    g545(.A(G50gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n721_), .B(new_n748_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n739_), .B2(new_n667_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT116), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n753_), .A3(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1331gat));
  NOR2_X1   g554(.A1(new_n697_), .A2(new_n492_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n681_), .A2(new_n638_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n582_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G57gat), .B1(new_n758_), .B2(new_n450_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT117), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n582_), .A2(new_n491_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n637_), .A2(new_n638_), .A3(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(G57gat), .A3(new_n450_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n760_), .A2(new_n763_), .ZN(G1332gat));
  INV_X1    g563(.A(G64gat), .ZN(new_n765_));
  INV_X1    g564(.A(new_n709_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n762_), .B2(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT48), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n758_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1333gat));
  INV_X1    g569(.A(G71gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n758_), .A2(new_n771_), .A3(new_n660_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n762_), .A2(new_n660_), .ZN(new_n773_));
  XOR2_X1   g572(.A(KEYINPUT118), .B(KEYINPUT49), .Z(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(G71gat), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G71gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  AOI21_X1  g576(.A(new_n548_), .B1(new_n762_), .B2(new_n668_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT50), .Z(new_n779_));
  NAND3_X1  g578(.A1(new_n758_), .A2(new_n548_), .A3(new_n668_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1335gat));
  NOR2_X1   g580(.A1(new_n761_), .A2(new_n624_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n364_), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n697_), .A2(new_n492_), .A3(new_n583_), .A4(new_n674_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n533_), .A3(new_n450_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1336gat));
  OAI21_X1  g586(.A(G92gat), .B1(new_n783_), .B2(new_n709_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n534_), .A3(new_n461_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n783_), .B2(new_n250_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n660_), .A3(new_n529_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n785_), .A2(new_n530_), .A3(new_n339_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n339_), .B(new_n782_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n796_));
  XOR2_X1   g595(.A(KEYINPUT119), .B(KEYINPUT52), .Z(new_n797_));
  AND3_X1   g596(.A1(new_n796_), .A2(G106gat), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n796_), .B2(G106gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n795_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  NOR2_X1   g603(.A1(new_n461_), .A2(new_n339_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n660_), .A3(new_n450_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n475_), .A2(new_n482_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n482_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n478_), .A2(new_n480_), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n811_), .A3(new_n488_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n490_), .A2(new_n812_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT120), .Z(new_n814_));
  INV_X1    g613(.A(new_n500_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n569_), .A2(new_n572_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n568_), .B1(new_n571_), .B2(KEYINPUT12), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n559_), .A2(new_n562_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n568_), .B(new_n559_), .C1(new_n571_), .C2(KEYINPUT12), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n561_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n558_), .A2(new_n563_), .A3(KEYINPUT55), .A4(new_n568_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n500_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n500_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n817_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n808_), .B1(new_n830_), .B2(KEYINPUT122), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n814_), .A2(new_n816_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n500_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n500_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n832_), .B(KEYINPUT122), .C1(new_n833_), .C2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n681_), .B1(new_n831_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT123), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n830_), .A2(KEYINPUT58), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n808_), .A3(new_n835_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n681_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n838_), .A2(new_n839_), .A3(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n816_), .A2(new_n492_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n578_), .A2(new_n814_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n673_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n850_), .A2(KEYINPUT57), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(KEYINPUT57), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n624_), .B1(new_n846_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT54), .B1(new_n625_), .B2(new_n492_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n757_), .A2(new_n857_), .A3(new_n491_), .A4(new_n583_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n807_), .B1(new_n855_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n845_), .A2(new_n839_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n844_), .B1(new_n843_), .B2(new_n681_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n852_), .A2(KEYINPUT121), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n851_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n850_), .A2(new_n867_), .A3(KEYINPUT57), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n638_), .B1(new_n864_), .B2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n806_), .B1(new_n871_), .B2(new_n859_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n492_), .B(new_n861_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G113gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n806_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n867_), .B1(new_n850_), .B2(KEYINPUT57), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n850_), .A2(KEYINPUT57), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n868_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n624_), .B1(new_n880_), .B2(new_n846_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n876_), .B1(new_n881_), .B2(new_n860_), .ZN(new_n882_));
  OR3_X1    g681(.A1(new_n882_), .A2(G113gat), .A3(new_n491_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n875_), .A2(new_n883_), .ZN(G1340gat));
  OAI211_X1 g683(.A(new_n582_), .B(new_n861_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G120gat), .ZN(new_n886_));
  INV_X1    g685(.A(G120gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n583_), .B2(KEYINPUT60), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT124), .B1(new_n887_), .B2(KEYINPUT60), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n872_), .B(new_n890_), .C1(new_n891_), .C2(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n886_), .A2(new_n892_), .ZN(G1341gat));
  OAI211_X1 g692(.A(new_n624_), .B(new_n861_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G127gat), .ZN(new_n895_));
  OR3_X1    g694(.A1(new_n882_), .A2(G127gat), .A3(new_n638_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1342gat));
  OAI211_X1 g696(.A(new_n673_), .B(new_n876_), .C1(new_n881_), .C2(new_n860_), .ZN(new_n898_));
  INV_X1    g697(.A(G134gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT125), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n898_), .A2(new_n902_), .A3(new_n899_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n846_), .A2(new_n854_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n638_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n859_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n882_), .A2(KEYINPUT59), .B1(new_n906_), .B2(new_n807_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n610_), .A2(new_n899_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n901_), .A2(new_n903_), .B1(new_n907_), .B2(new_n908_), .ZN(G1343gat));
  NAND2_X1  g708(.A1(new_n871_), .A2(new_n859_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n766_), .A2(new_n660_), .A3(new_n746_), .A4(new_n364_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n492_), .A3(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n582_), .A3(new_n911_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n910_), .A2(new_n624_), .A3(new_n911_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n911_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G162gat), .B1(new_n919_), .B2(new_n610_), .ZN(new_n920_));
  INV_X1    g719(.A(G162gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n673_), .A2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n919_), .B2(new_n922_), .ZN(G1347gat));
  NOR3_X1   g722(.A1(new_n709_), .A2(new_n250_), .A3(new_n450_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n668_), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n492_), .B(new_n926_), .C1(new_n855_), .C2(new_n860_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n221_), .B1(new_n928_), .B2(KEYINPUT62), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(KEYINPUT126), .A3(new_n931_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n927_), .B(new_n929_), .C1(new_n928_), .C2(KEYINPUT62), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n932_), .B(new_n933_), .C1(new_n374_), .C2(new_n927_), .ZN(G1348gat));
  NOR2_X1   g733(.A1(new_n855_), .A2(new_n860_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n926_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G176gat), .B1(new_n937_), .B2(new_n582_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n881_), .A2(new_n860_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n339_), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n924_), .A2(G176gat), .A3(new_n582_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n938_), .B1(new_n940_), .B2(new_n941_), .ZN(G1349gat));
  NAND3_X1  g741(.A1(new_n940_), .A2(new_n624_), .A3(new_n924_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n638_), .A2(new_n212_), .ZN(new_n944_));
  AOI22_X1  g743(.A1(new_n943_), .A2(new_n377_), .B1(new_n937_), .B2(new_n944_), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n937_), .A2(new_n213_), .A3(new_n673_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n935_), .A2(new_n610_), .A3(new_n936_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n381_), .ZN(G1351gat));
  NOR3_X1   g747(.A1(new_n746_), .A2(new_n660_), .A3(new_n450_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n766_), .A2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n939_), .A2(new_n950_), .ZN(new_n951_));
  AND3_X1   g750(.A1(new_n951_), .A2(G197gat), .A3(new_n492_), .ZN(new_n952_));
  AOI21_X1  g751(.A(G197gat), .B1(new_n951_), .B2(new_n492_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1352gat));
  NAND3_X1  g753(.A1(new_n910_), .A2(new_n766_), .A3(new_n949_), .ZN(new_n955_));
  OAI21_X1  g754(.A(G204gat), .B1(new_n955_), .B2(new_n583_), .ZN(new_n956_));
  INV_X1    g755(.A(G204gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n951_), .A2(new_n957_), .A3(new_n582_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n956_), .A2(new_n958_), .ZN(G1353gat));
  NOR3_X1   g758(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960_));
  AOI211_X1 g759(.A(new_n960_), .B(new_n638_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n951_), .A2(new_n961_), .ZN(new_n962_));
  OAI21_X1  g761(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n951_), .A2(new_n963_), .A3(new_n961_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1354gat));
  OAI21_X1  g766(.A(G218gat), .B1(new_n955_), .B2(new_n610_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n951_), .A2(new_n264_), .A3(new_n673_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1355gat));
endmodule


