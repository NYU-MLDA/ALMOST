//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n985_, new_n986_, new_n987_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n995_, new_n996_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1003_, new_n1004_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT19), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G211gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G218gat), .ZN(new_n210_));
  INV_X1    g009(.A(G218gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(G211gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT85), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G197gat), .A2(G204gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G197gat), .A2(G204gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(G211gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n209_), .A2(G218gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT85), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n213_), .A2(new_n218_), .A3(new_n222_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n221_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n216_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(KEYINPUT21), .A3(new_n214_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n217_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n223_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT86), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT23), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(G183gat), .A3(G190gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n235_), .A2(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT76), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G169gat), .A3(G176gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n242_), .A2(new_n244_), .A3(new_n245_), .A4(KEYINPUT24), .ZN(new_n246_));
  INV_X1    g045(.A(G183gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT25), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G183gat), .ZN(new_n250_));
  INV_X1    g049(.A(G190gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT26), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT26), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G190gat), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n248_), .A2(new_n250_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n240_), .A2(new_n246_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT77), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT22), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(G169gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT22), .B(G169gat), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n257_), .B(new_n260_), .C1(new_n261_), .C2(new_n258_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n243_), .B1(G169gat), .B2(G176gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n241_), .A2(KEYINPUT76), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n235_), .A2(new_n237_), .A3(KEYINPUT78), .ZN(new_n267_));
  OR3_X1    g066(.A1(new_n234_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n247_), .A2(new_n251_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n256_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n228_), .B(new_n229_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT86), .A3(new_n223_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n233_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n272_), .A2(KEYINPUT87), .A3(new_n223_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT87), .B1(new_n272_), .B2(new_n223_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n238_), .A2(KEYINPUT89), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT89), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT24), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n282_), .A3(new_n239_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n255_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n267_), .A2(new_n268_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n245_), .A2(new_n241_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n284_), .A2(new_n285_), .A3(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT90), .B1(new_n263_), .B2(new_n264_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n242_), .A2(new_n244_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n235_), .A2(new_n237_), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n294_), .A2(new_n269_), .B1(new_n261_), .B2(new_n257_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n289_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n276_), .B1(new_n279_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT95), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n275_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n231_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n272_), .A2(KEYINPUT87), .A3(new_n223_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n284_), .A2(new_n288_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n285_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n236_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n234_), .A2(KEYINPUT23), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n269_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n261_), .A2(new_n257_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n242_), .A2(new_n244_), .A3(new_n291_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n291_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n309_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n301_), .A2(new_n302_), .A3(new_n305_), .A4(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT20), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT95), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n208_), .B1(new_n299_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n233_), .A2(new_n273_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n271_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n276_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n293_), .A2(new_n320_), .A3(new_n295_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n305_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT92), .A3(new_n231_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n312_), .A2(KEYINPUT91), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n293_), .A2(new_n320_), .A3(new_n295_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n289_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n272_), .A2(new_n223_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n325_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AND4_X1   g129(.A1(new_n208_), .A2(new_n319_), .A3(new_n324_), .A4(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n205_), .B1(new_n316_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT27), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n329_), .B(new_n305_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n207_), .A2(new_n276_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n274_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n319_), .A2(new_n330_), .A3(new_n324_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n207_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n205_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n333_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n332_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n207_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n336_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n339_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  AOI211_X1 g143(.A(new_n205_), .B(new_n336_), .C1(new_n337_), .C2(new_n207_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n333_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G78gat), .B(G106gat), .Z(new_n347_));
  AND2_X1   g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT2), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(KEYINPUT2), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n355_), .A2(new_n351_), .B1(G141gat), .B2(G148gat), .ZN(new_n356_));
  OR2_X1    g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357_));
  OAI22_X1  g156(.A1(new_n354_), .A2(new_n356_), .B1(KEYINPUT3), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n350_), .A2(KEYINPUT3), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n348_), .A2(new_n349_), .A3(KEYINPUT1), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT82), .ZN(new_n362_));
  NAND3_X1  g161(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n352_), .A3(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n359_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n350_), .A2(new_n358_), .B1(new_n365_), .B2(new_n357_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n357_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n353_), .B1(new_n361_), .B2(KEYINPUT82), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n351_), .B1(new_n372_), .B2(KEYINPUT83), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n371_), .A2(new_n372_), .B1(new_n373_), .B2(new_n361_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n357_), .A2(KEYINPUT3), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n350_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n370_), .A2(new_n368_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT28), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n369_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n369_), .B2(new_n378_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n370_), .A2(new_n376_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT29), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n278_), .B2(new_n277_), .ZN(new_n386_));
  INV_X1    g185(.A(G233gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n387_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n233_), .A2(new_n393_), .A3(new_n273_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n385_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n347_), .B1(new_n383_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n383_), .A2(new_n396_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n369_), .A2(new_n378_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n379_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n380_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n386_), .A2(new_n391_), .B1(new_n394_), .B2(new_n385_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n347_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .A4(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n398_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n406_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n405_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n341_), .A2(new_n346_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G85gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT0), .B(G57gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n414_), .B(new_n415_), .Z(new_n416_));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G127gat), .B(G134gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G113gat), .B(G120gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT81), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n418_), .B(new_n419_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT81), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n384_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n370_), .A2(new_n422_), .A3(new_n376_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n417_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT4), .B1(new_n384_), .B2(new_n424_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n428_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n416_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n418_), .A2(new_n419_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n418_), .A2(new_n419_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n423_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n420_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n426_), .B1(new_n366_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT4), .ZN(new_n439_));
  INV_X1    g238(.A(new_n429_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n431_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n416_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n432_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n433_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n318_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n271_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT80), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n424_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(KEYINPUT80), .A3(new_n437_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT80), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n447_), .A2(new_n455_), .A3(new_n449_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457_));
  INV_X1    g256(.A(G43gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G227gat), .A2(G233gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(G15gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n459_), .B(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT31), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT31), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n466_), .A3(new_n462_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n454_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n464_), .A2(new_n452_), .A3(new_n467_), .A4(new_n453_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n445_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT98), .B1(new_n412_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n342_), .A2(new_n343_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n205_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n338_), .A2(new_n339_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n476_), .A2(new_n333_), .B1(new_n332_), .B2(new_n340_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n409_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n397_), .A2(new_n406_), .B1(new_n399_), .B2(new_n398_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n471_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT98), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n477_), .A2(new_n480_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n472_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n474_), .A2(new_n485_), .A3(new_n475_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT93), .B1(new_n344_), .B2(new_n345_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n442_), .B1(new_n438_), .B2(new_n428_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n429_), .B1(new_n438_), .B2(KEYINPUT4), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n488_), .B1(new_n490_), .B2(new_n428_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n432_), .B1(new_n489_), .B2(new_n431_), .ZN(new_n492_));
  OAI22_X1  g291(.A1(new_n492_), .A2(new_n442_), .B1(KEYINPUT94), .B2(KEYINPUT33), .ZN(new_n493_));
  NOR2_X1   g292(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n416_), .B(new_n494_), .C1(new_n430_), .C2(new_n432_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n491_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n486_), .A2(new_n487_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n339_), .A2(KEYINPUT32), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n338_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n433_), .A2(new_n444_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n313_), .A2(new_n298_), .A3(KEYINPUT20), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n315_), .A2(new_n274_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n331_), .B1(new_n207_), .B2(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n499_), .B(new_n500_), .C1(new_n503_), .C2(new_n498_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT32), .B(new_n339_), .C1(new_n316_), .C2(new_n331_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n507_), .A2(KEYINPUT96), .A3(new_n499_), .A4(new_n500_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n497_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n480_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n445_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n341_), .A2(new_n346_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT97), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n500_), .B1(new_n411_), .B2(new_n407_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT97), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n477_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n510_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n469_), .A2(new_n470_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n484_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G29gat), .B(G36gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT71), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT71), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT15), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530_));
  INV_X1    g329(.A(G1gat), .ZN(new_n531_));
  INV_X1    g330(.A(G8gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT14), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G8gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n529_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n528_), .B2(new_n536_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n528_), .B(new_n537_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(new_n539_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OR3_X1    g346(.A1(new_n541_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n519_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n556_));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT64), .B(G85gat), .Z(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT9), .B1(new_n566_), .B2(G92gat), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n567_), .B2(KEYINPUT65), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT64), .B(G85gat), .ZN(new_n569_));
  INV_X1    g368(.A(G92gat), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n563_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT65), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT6), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(G106gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT10), .B(G99gat), .Z(new_n579_));
  AOI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n577_), .B1(KEYINPUT66), .B2(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(KEYINPUT66), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n562_), .A2(new_n564_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT8), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n562_), .B(new_n564_), .C1(new_n577_), .C2(new_n586_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n589_), .A2(new_n592_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n560_), .B1(new_n581_), .B2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n581_), .A2(new_n594_), .A3(new_n560_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT67), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT67), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n581_), .A2(new_n594_), .A3(new_n598_), .A4(new_n560_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n595_), .B1(new_n600_), .B2(KEYINPUT68), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT68), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n602_), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n595_), .A2(KEYINPUT12), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT69), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n591_), .B(new_n590_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n593_), .A2(new_n591_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n594_), .A2(KEYINPUT69), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n581_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n560_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT12), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n608_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n605_), .A3(new_n596_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT5), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n607_), .A2(new_n620_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n605_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n612_), .A2(new_n613_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n628_));
  OAI22_X1  g427(.A1(new_n628_), .A2(new_n617_), .B1(KEYINPUT12), .B2(new_n595_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n596_), .A2(new_n605_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n624_), .B1(new_n627_), .B2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n632_), .A3(KEYINPUT70), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT70), .B1(new_n626_), .B2(new_n632_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n553_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT70), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n625_), .B1(new_n607_), .B2(new_n620_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n627_), .A2(new_n631_), .A3(new_n624_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(KEYINPUT13), .A3(new_n633_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT34), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT72), .B1(new_n644_), .B2(KEYINPUT35), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n581_), .A2(new_n594_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n528_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n648_), .B1(new_n529_), .B2(new_n628_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n644_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT35), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n652_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n648_), .B(new_n654_), .C1(new_n529_), .C2(new_n628_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G190gat), .B(G218gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT36), .Z(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT74), .Z(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT75), .B1(new_n656_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT75), .ZN(new_n664_));
  AOI211_X1 g463(.A(new_n664_), .B(new_n661_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n659_), .A2(KEYINPUT36), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n653_), .A2(new_n667_), .A3(new_n655_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT73), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT73), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n653_), .A2(new_n670_), .A3(new_n667_), .A4(new_n655_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT37), .B1(new_n666_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT37), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n656_), .B2(new_n662_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n672_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n537_), .B(new_n560_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(G231gat), .A2(G233gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT17), .ZN(new_n681_));
  XOR2_X1   g480(.A(G127gat), .B(G155gat), .Z(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT16), .ZN(new_n683_));
  XNOR2_X1  g482(.A(G183gat), .B(G211gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n680_), .A2(new_n681_), .A3(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(KEYINPUT17), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n680_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n673_), .A2(new_n676_), .A3(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n552_), .A2(new_n642_), .A3(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n691_), .A2(G1gat), .A3(new_n445_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n692_), .A2(KEYINPUT38), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(KEYINPUT38), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n656_), .A2(new_n662_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n664_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n656_), .A2(KEYINPUT75), .A3(new_n662_), .ZN(new_n697_));
  AND4_X1   g496(.A1(KEYINPUT99), .A2(new_n672_), .A3(new_n696_), .A4(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT99), .B1(new_n666_), .B2(new_n672_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n519_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n689_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n702_), .A2(new_n550_), .A3(new_n642_), .A4(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G1gat), .B1(new_n704_), .B2(new_n445_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n693_), .A2(new_n694_), .A3(new_n705_), .ZN(G1324gat));
  NOR3_X1   g505(.A1(new_n691_), .A2(G8gat), .A3(new_n477_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G8gat), .B1(new_n704_), .B2(new_n477_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n708_), .A2(KEYINPUT39), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(KEYINPUT39), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n711_), .B(new_n712_), .Z(G1325gat));
  OAI21_X1  g512(.A(G15gat), .B1(new_n704_), .B2(new_n518_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT41), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n691_), .A2(G15gat), .A3(new_n518_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1326gat));
  XOR2_X1   g516(.A(new_n480_), .B(KEYINPUT101), .Z(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G22gat), .B1(new_n704_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT42), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n719_), .A2(G22gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n691_), .B2(new_n722_), .ZN(G1327gat));
  NAND3_X1  g522(.A1(new_n642_), .A2(new_n550_), .A3(new_n689_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n509_), .A2(new_n480_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n513_), .A2(new_n516_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n518_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n484_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n672_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n733_), .A2(new_n674_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n727_), .B1(new_n732_), .B2(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n519_), .A2(KEYINPUT43), .A3(new_n734_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n725_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n726_), .B1(new_n519_), .B2(new_n734_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n743_));
  INV_X1    g542(.A(new_n518_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n513_), .A2(new_n516_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n510_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n743_), .B(new_n735_), .C1(new_n746_), .C2(new_n484_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n724_), .B1(new_n742_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT103), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n740_), .A2(new_n741_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(KEYINPUT44), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752_), .B2(new_n445_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT104), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT104), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n700_), .A2(new_n703_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n642_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n552_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n445_), .A2(G29gat), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n754_), .A2(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1328gat));
  NAND2_X1  g559(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT108), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n477_), .B1(new_n748_), .B2(KEYINPUT44), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n741_), .B1(new_n748_), .B2(KEYINPUT103), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n739_), .B(new_n724_), .C1(new_n742_), .C2(new_n747_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT105), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n766_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(G36gat), .A3(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n477_), .A2(G36gat), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT106), .B1(new_n758_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n757_), .A2(new_n552_), .A3(new_n777_), .A4(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT45), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n762_), .B(new_n765_), .C1(new_n773_), .C2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n772_), .A2(G36gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n771_), .B1(new_n750_), .B2(new_n766_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n764_), .B1(new_n784_), .B2(new_n761_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n781_), .A2(new_n785_), .ZN(G1329gat));
  OAI21_X1  g585(.A(new_n458_), .B1(new_n758_), .B2(new_n518_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n744_), .A2(G43gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n752_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g589(.A(G50gat), .B1(new_n752_), .B2(new_n480_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n719_), .A2(G50gat), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT109), .Z(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n758_), .B2(new_n793_), .ZN(G1331gat));
  NOR3_X1   g593(.A1(new_n642_), .A2(new_n550_), .A3(new_n689_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n702_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT110), .B(G57gat), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n445_), .A3(new_n797_), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT111), .Z(new_n799_));
  NOR2_X1   g598(.A1(new_n642_), .A2(new_n550_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n732_), .A2(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n801_), .A2(new_n689_), .A3(new_n735_), .ZN(new_n802_));
  AOI21_X1  g601(.A(G57gat), .B1(new_n802_), .B2(new_n500_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n799_), .A2(new_n803_), .ZN(G1332gat));
  OAI21_X1  g603(.A(G64gat), .B1(new_n796_), .B2(new_n477_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT48), .ZN(new_n806_));
  INV_X1    g605(.A(G64gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n802_), .A2(new_n807_), .A3(new_n512_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1333gat));
  OAI21_X1  g608(.A(G71gat), .B1(new_n796_), .B2(new_n518_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT49), .ZN(new_n811_));
  INV_X1    g610(.A(G71gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n802_), .A2(new_n812_), .A3(new_n744_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1334gat));
  INV_X1    g613(.A(G78gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n802_), .A2(new_n815_), .A3(new_n718_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n702_), .A2(new_n718_), .A3(new_n795_), .ZN(new_n817_));
  XOR2_X1   g616(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n818_));
  AND3_X1   g617(.A1(new_n817_), .A2(G78gat), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n817_), .B2(G78gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(G1335gat));
  INV_X1    g620(.A(new_n801_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n756_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G85gat), .B1(new_n824_), .B2(new_n500_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n551_), .A2(new_n689_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n642_), .B(new_n826_), .C1(new_n742_), .C2(new_n747_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n445_), .A2(new_n569_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n825_), .B1(new_n827_), .B2(new_n828_), .ZN(G1336gat));
  NAND3_X1  g628(.A1(new_n824_), .A2(new_n570_), .A3(new_n512_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n827_), .A2(new_n512_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n570_), .ZN(G1337gat));
  INV_X1    g631(.A(G99gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n827_), .B2(new_n744_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n824_), .A2(new_n744_), .A3(new_n579_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n836_));
  OAI22_X1  g635(.A1(new_n834_), .A2(new_n835_), .B1(new_n836_), .B2(KEYINPUT51), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(KEYINPUT51), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1338gat));
  INV_X1    g638(.A(new_n480_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n824_), .A2(new_n578_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n827_), .A2(new_n840_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(G106gat), .ZN(new_n844_));
  AOI211_X1 g643(.A(KEYINPUT52), .B(new_n578_), .C1(new_n827_), .C2(new_n840_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n550_), .A2(G113gat), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT120), .Z(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n642_), .A2(new_n690_), .A3(new_n551_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n852_), .A2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n853_), .B(KEYINPUT115), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n642_), .A2(new_n690_), .A3(new_n551_), .A4(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n626_), .A2(new_n550_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n619_), .A2(KEYINPUT117), .A3(new_n597_), .A4(new_n599_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n629_), .B2(new_n600_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n863_), .A3(new_n606_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT55), .B1(new_n631_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n620_), .A2(KEYINPUT116), .A3(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n866_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n624_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(KEYINPUT56), .A3(new_n624_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n860_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n539_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n528_), .B2(new_n536_), .ZN(new_n876_));
  OAI221_X1 g675(.A(new_n547_), .B1(new_n542_), .B2(new_n875_), .C1(new_n538_), .C2(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n548_), .A2(new_n877_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n640_), .A2(new_n633_), .A3(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n700_), .B1(new_n874_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n700_), .B(KEYINPUT57), .C1(new_n874_), .C2(new_n879_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n878_), .A2(new_n626_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n869_), .A2(KEYINPUT56), .A3(new_n624_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n869_), .B2(new_n624_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT58), .B(new_n884_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n735_), .A3(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n882_), .A2(new_n883_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n859_), .B1(new_n689_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n412_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n518_), .A2(new_n445_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n896_), .A2(KEYINPUT119), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(KEYINPUT119), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n893_), .A2(KEYINPUT59), .A3(new_n897_), .A4(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n893_), .A2(new_n896_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT118), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n903_), .B(KEYINPUT59), .C1(new_n893_), .C2(new_n896_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n851_), .B(new_n899_), .C1(new_n902_), .C2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G113gat), .B1(new_n900_), .B2(new_n550_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n848_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n899_), .B1(new_n902_), .B2(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n850_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n906_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(KEYINPUT121), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n907_), .A2(new_n911_), .ZN(G1340gat));
  INV_X1    g711(.A(G120gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n642_), .B2(KEYINPUT60), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n900_), .B(new_n914_), .C1(KEYINPUT60), .C2(new_n913_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n642_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n908_), .A2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n917_), .B2(new_n913_), .ZN(G1341gat));
  INV_X1    g717(.A(G127gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n900_), .A2(new_n919_), .A3(new_n703_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n908_), .A2(new_n703_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n919_), .ZN(G1342gat));
  INV_X1    g721(.A(G134gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n900_), .A2(new_n923_), .A3(new_n701_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n908_), .A2(new_n735_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(G1343gat));
  NOR2_X1   g725(.A1(new_n480_), .A2(new_n744_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n512_), .A2(new_n445_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n734_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n929_));
  AOI22_X1  g728(.A1(new_n881_), .A2(new_n880_), .B1(new_n929_), .B2(new_n890_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n703_), .B1(new_n930_), .B2(new_n883_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n927_), .B(new_n928_), .C1(new_n931_), .C2(new_n859_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n892_), .A2(new_n689_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n859_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n937_), .A2(KEYINPUT122), .A3(new_n927_), .A4(new_n928_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n934_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n550_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n916_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g742(.A(new_n938_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n927_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n945_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n946_));
  AOI21_X1  g745(.A(KEYINPUT122), .B1(new_n946_), .B2(new_n928_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n703_), .B1(new_n944_), .B2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(KEYINPUT123), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n939_), .A2(new_n950_), .A3(new_n703_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT61), .B(G155gat), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n949_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n952_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n950_), .B1(new_n939_), .B2(new_n703_), .ZN(new_n955_));
  AOI211_X1 g754(.A(KEYINPUT123), .B(new_n689_), .C1(new_n934_), .C2(new_n938_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n954_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n953_), .A2(new_n957_), .ZN(G1346gat));
  INV_X1    g757(.A(new_n939_), .ZN(new_n959_));
  OR3_X1    g758(.A1(new_n959_), .A2(G162gat), .A3(new_n700_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G162gat), .B1(new_n959_), .B2(new_n734_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1347gat));
  NOR2_X1   g761(.A1(new_n477_), .A2(new_n500_), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n718_), .A2(new_n518_), .A3(new_n964_), .ZN(new_n965_));
  AND2_X1   g764(.A1(new_n937_), .A2(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n550_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n967_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n968_));
  INV_X1    g767(.A(new_n261_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n968_), .B1(new_n969_), .B2(new_n967_), .ZN(new_n970_));
  AOI21_X1  g769(.A(KEYINPUT62), .B1(new_n967_), .B2(G169gat), .ZN(new_n971_));
  OR2_X1    g770(.A1(new_n970_), .A2(new_n971_), .ZN(G1348gat));
  AOI21_X1  g771(.A(G176gat), .B1(new_n966_), .B2(new_n916_), .ZN(new_n973_));
  AOI21_X1  g772(.A(KEYINPUT124), .B1(new_n937_), .B2(new_n480_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n975_));
  NOR3_X1   g774(.A1(new_n893_), .A2(new_n975_), .A3(new_n840_), .ZN(new_n976_));
  NOR4_X1   g775(.A1(new_n974_), .A2(new_n976_), .A3(new_n518_), .A4(new_n964_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n642_), .A2(new_n257_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n973_), .B1(new_n977_), .B2(new_n978_), .ZN(G1349gat));
  AOI21_X1  g778(.A(new_n689_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n966_), .A2(new_n980_), .ZN(new_n981_));
  XOR2_X1   g780(.A(new_n981_), .B(KEYINPUT125), .Z(new_n982_));
  AOI21_X1  g781(.A(G183gat), .B1(new_n977_), .B2(new_n703_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n982_), .A2(new_n983_), .ZN(G1350gat));
  INV_X1    g783(.A(new_n966_), .ZN(new_n985_));
  OAI21_X1  g784(.A(G190gat), .B1(new_n985_), .B2(new_n734_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n701_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n986_), .B1(new_n985_), .B2(new_n987_), .ZN(G1351gat));
  XNOR2_X1  g787(.A(KEYINPUT126), .B(G197gat), .ZN(new_n989_));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n990_), .A2(G197gat), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n946_), .A2(new_n963_), .ZN(new_n992_));
  NOR2_X1   g791(.A1(new_n992_), .A2(new_n551_), .ZN(new_n993_));
  MUX2_X1   g792(.A(new_n989_), .B(new_n991_), .S(new_n993_), .Z(G1352gat));
  INV_X1    g793(.A(new_n992_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n995_), .A2(new_n916_), .ZN(new_n996_));
  XNOR2_X1  g795(.A(new_n996_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g796(.A1(new_n992_), .A2(new_n689_), .ZN(new_n998_));
  NOR2_X1   g797(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n999_));
  AND2_X1   g798(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1000_));
  OAI21_X1  g799(.A(new_n998_), .B1(new_n999_), .B2(new_n1000_), .ZN(new_n1001_));
  OAI21_X1  g800(.A(new_n1001_), .B1(new_n998_), .B2(new_n999_), .ZN(G1354gat));
  OAI21_X1  g801(.A(G218gat), .B1(new_n992_), .B2(new_n734_), .ZN(new_n1003_));
  NAND2_X1  g802(.A1(new_n701_), .A2(new_n211_), .ZN(new_n1004_));
  OAI21_X1  g803(.A(new_n1003_), .B1(new_n992_), .B2(new_n1004_), .ZN(G1355gat));
endmodule


