//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_;
  XNOR2_X1  g000(.A(KEYINPUT69), .B(G71gat), .ZN(new_n202_));
  INV_X1    g001(.A(G78gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(KEYINPUT11), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT70), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G85gat), .B(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n217_), .C1(G99gat), .C2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n219_), .B(new_n220_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT68), .Z(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT6), .B1(new_n219_), .B2(new_n220_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT6), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT67), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n215_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n213_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT71), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT9), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G85gat), .A3(G92gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n227_), .B(new_n236_), .C1(new_n235_), .C2(new_n213_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT10), .B(G99gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT65), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n239_), .B2(new_n220_), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT72), .Z(new_n241_));
  NAND2_X1  g040(.A1(new_n234_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n232_), .A2(new_n233_), .ZN(new_n243_));
  OAI211_X1 g042(.A(KEYINPUT12), .B(new_n212_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n239_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G106gat), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n229_), .B(new_n231_), .C1(new_n246_), .C2(new_n237_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT12), .B1(new_n212_), .B2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n212_), .A2(new_n247_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT64), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n244_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n252_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n247_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(new_n211_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n256_), .B2(new_n249_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G120gat), .B(G148gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT5), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G176gat), .B(G204gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(new_n257_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT13), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(KEYINPUT13), .A3(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271_));
  INV_X1    g070(.A(G1gat), .ZN(new_n272_));
  INV_X1    g071(.A(G8gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT14), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G1gat), .B(G8gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G29gat), .B(G36gat), .Z(new_n279_));
  XOR2_X1   g078(.A(G43gat), .B(G50gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n281_), .B(KEYINPUT15), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(new_n277_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G229gat), .A2(G233gat), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n281_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n277_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n288_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G113gat), .B(G141gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G169gat), .B(G197gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT77), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n294_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n270_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n306_));
  NOR2_X1   g105(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G183gat), .ZN(new_n309_));
  INV_X1    g108(.A(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n311_), .C1(KEYINPUT23), .C2(new_n305_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT22), .B(G169gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT79), .ZN(new_n316_));
  INV_X1    g115(.A(G176gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n317_), .B1(new_n316_), .B2(KEYINPUT22), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G169gat), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n323_), .B2(new_n305_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(KEYINPUT80), .A3(new_n311_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n314_), .A2(new_n321_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n304_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n305_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT25), .B(G183gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G190gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n331_), .A2(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT24), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n330_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n326_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G227gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G15gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n340_), .B(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G127gat), .B(G134gat), .Z(new_n344_));
  XOR2_X1   g143(.A(G113gat), .B(G120gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n343_), .B(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G71gat), .B(G99gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT82), .B(G43gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n347_), .B(new_n354_), .Z(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT91), .Z(new_n358_));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT85), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n361_));
  INV_X1    g160(.A(G141gat), .ZN(new_n362_));
  INV_X1    g161(.A(G148gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n360_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n367_), .A2(KEYINPUT84), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(KEYINPUT84), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT85), .B(new_n366_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G141gat), .A2(G148gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT2), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(G141gat), .A3(G148gat), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n372_), .A2(new_n374_), .B1(new_n364_), .B2(KEYINPUT3), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n365_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n378_), .A2(KEYINPUT86), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT86), .B1(new_n378_), .B2(new_n379_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n377_), .B1(KEYINPUT1), .B2(new_n379_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n384_), .B1(KEYINPUT1), .B2(new_n379_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n364_), .A3(new_n371_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n383_), .A2(KEYINPUT87), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT87), .B1(new_n383_), .B2(new_n386_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n359_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT28), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT28), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n391_), .B(new_n359_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n358_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n392_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n393_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n358_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n383_), .A2(new_n386_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT87), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n383_), .A2(KEYINPUT87), .A3(new_n386_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT29), .A3(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G211gat), .B(G218gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(G197gat), .A2(G204gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G197gat), .A2(G204gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(KEYINPUT21), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT21), .B1(new_n411_), .B2(new_n412_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G211gat), .B(G218gat), .Z(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n410_), .B(new_n413_), .C1(new_n416_), .C2(new_n415_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n418_), .A2(KEYINPUT90), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT90), .B1(new_n418_), .B2(new_n419_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n407_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT88), .Z(new_n425_));
  AND2_X1   g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n418_), .A2(new_n419_), .ZN(new_n427_));
  AOI211_X1 g226(.A(new_n425_), .B(new_n427_), .C1(new_n403_), .C2(KEYINPUT29), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n396_), .A2(new_n402_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n396_), .B2(new_n402_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n331_), .A2(new_n332_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n334_), .A2(new_n333_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n338_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n324_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT92), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT92), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n335_), .A2(new_n438_), .A3(new_n324_), .A4(new_n338_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT93), .ZN(new_n441_));
  INV_X1    g240(.A(new_n311_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n315_), .A2(new_n317_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n337_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n441_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n330_), .A2(new_n311_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n445_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(KEYINPUT93), .A3(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n440_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n427_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G226gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT19), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n339_), .B(new_n326_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n452_), .A2(KEYINPUT20), .A3(new_n455_), .A4(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT99), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n422_), .B2(new_n340_), .ZN(new_n461_));
  OAI221_X1 g260(.A(new_n427_), .B1(new_n435_), .B2(new_n436_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n454_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n427_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n418_), .A2(KEYINPUT90), .A3(new_n419_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n326_), .A2(new_n339_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n460_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(KEYINPUT99), .A3(new_n452_), .A4(new_n455_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n459_), .A2(new_n464_), .A3(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G8gat), .B(G36gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(G64gat), .B(G92gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n477_), .A2(KEYINPUT32), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n455_), .B1(new_n470_), .B2(new_n452_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n340_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n440_), .A2(new_n427_), .A3(new_n446_), .A4(new_n449_), .ZN(new_n482_));
  AND4_X1   g281(.A1(KEYINPUT20), .A2(new_n481_), .A3(new_n482_), .A4(new_n455_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n479_), .B1(new_n485_), .B2(new_n478_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G1gat), .B(G29gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G57gat), .B(G85gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  NAND2_X1  g290(.A1(G225gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n346_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n405_), .A2(new_n493_), .A3(new_n406_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(KEYINPUT4), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n383_), .A2(new_n346_), .A3(new_n386_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT95), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n383_), .A2(new_n498_), .A3(new_n346_), .A4(new_n386_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n494_), .A2(new_n500_), .A3(KEYINPUT4), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n495_), .B1(new_n501_), .B2(KEYINPUT96), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT96), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n494_), .A2(new_n500_), .A3(new_n503_), .A4(KEYINPUT4), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n492_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n494_), .A2(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n492_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n491_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n501_), .A2(KEYINPUT96), .ZN(new_n510_));
  INV_X1    g309(.A(new_n495_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n504_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n508_), .B1(new_n512_), .B2(new_n507_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n491_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n486_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT33), .B1(new_n513_), .B2(new_n514_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT33), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n518_), .B(new_n491_), .C1(new_n505_), .C2(new_n508_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n491_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n512_), .B2(new_n507_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n477_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n456_), .A2(KEYINPUT20), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n449_), .A2(new_n446_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n427_), .B1(new_n526_), .B2(new_n440_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n454_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n461_), .A2(new_n455_), .A3(new_n482_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n477_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n522_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n520_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n516_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n532_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT98), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n432_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n472_), .A2(new_n523_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT27), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n484_), .B2(new_n477_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n524_), .A2(new_n530_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n540_), .A2(new_n542_), .B1(new_n543_), .B2(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n396_), .A2(new_n402_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n429_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n396_), .A2(new_n402_), .A3(new_n429_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n515_), .A2(new_n509_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT100), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n515_), .A2(new_n509_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT100), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n552_), .A2(new_n432_), .A3(new_n553_), .A4(new_n544_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n356_), .B1(new_n539_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n548_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n355_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n544_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(new_n550_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n303_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n284_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT34), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT35), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n255_), .A2(new_n281_), .B1(new_n568_), .B2(new_n567_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n570_), .B1(new_n564_), .B2(new_n571_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT73), .ZN(new_n576_));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT36), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n578_), .A2(new_n579_), .ZN(new_n582_));
  OAI22_X1  g381(.A1(new_n573_), .A2(new_n574_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n574_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n580_), .A3(new_n572_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n586_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT37), .B1(new_n586_), .B2(KEYINPUT74), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n277_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n211_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT16), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT17), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  OR3_X1    g400(.A1(new_n594_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NOR4_X1   g401(.A1(new_n593_), .A2(KEYINPUT75), .A3(new_n599_), .A4(new_n598_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT75), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n594_), .B2(new_n600_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n602_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n590_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n563_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n550_), .A2(new_n272_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n608_), .A2(KEYINPUT101), .A3(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT101), .B1(new_n608_), .B2(new_n609_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT38), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n586_), .A2(new_n606_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n486_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n550_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n537_), .B2(KEYINPUT98), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n535_), .B(new_n532_), .C1(new_n517_), .C2(new_n519_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n557_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n551_), .A2(new_n554_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n355_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n302_), .B(new_n614_), .C1(new_n621_), .C2(new_n561_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n552_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n612_), .A2(KEYINPUT38), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n613_), .A2(new_n627_), .A3(new_n628_), .ZN(G1324gat));
  OAI21_X1  g428(.A(G8gat), .B1(new_n622_), .B2(new_n544_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n608_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n544_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n273_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n636_), .B(new_n638_), .ZN(G1325gat));
  OAI21_X1  g438(.A(G15gat), .B1(new_n626_), .B2(new_n356_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n608_), .A2(G15gat), .A3(new_n356_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1326gat));
  INV_X1    g443(.A(G22gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n432_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT106), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n633_), .A2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n649_));
  OAI21_X1  g448(.A(new_n432_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(G22gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n534_), .A2(new_n535_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n538_), .A3(new_n616_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n555_), .B1(new_n653_), .B2(new_n557_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n562_), .B1(new_n654_), .B2(new_n355_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n655_), .A2(KEYINPUT102), .A3(new_n302_), .A4(new_n614_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n622_), .A2(new_n623_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n557_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n649_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n658_), .A2(new_n645_), .A3(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n648_), .B1(new_n651_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT107), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n648_), .B(new_n663_), .C1(new_n651_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1327gat));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  INV_X1    g465(.A(new_n588_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n586_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT108), .B1(new_n587_), .B2(new_n588_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(new_n621_), .B2(new_n561_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n589_), .A2(KEYINPUT43), .ZN(new_n674_));
  AOI22_X1  g473(.A1(KEYINPUT43), .A2(new_n673_), .B1(new_n655_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n606_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n303_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n666_), .B1(new_n675_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n655_), .B2(new_n672_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n621_), .A2(new_n561_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n674_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT44), .B(new_n677_), .C1(new_n681_), .C2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n679_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(G29gat), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n552_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n586_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n676_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n563_), .A2(new_n550_), .A3(new_n690_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n686_), .A2(new_n688_), .B1(new_n687_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(KEYINPUT109), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n679_), .A2(new_n634_), .A3(new_n685_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n544_), .A2(G36gat), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n563_), .A2(new_n698_), .A3(new_n690_), .A4(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n302_), .B(new_n690_), .C1(new_n621_), .C2(new_n561_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n699_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT45), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n693_), .A2(KEYINPUT109), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n695_), .B1(new_n697_), .B2(new_n707_), .ZN(new_n708_));
  AOI211_X1 g507(.A(new_n694_), .B(new_n706_), .C1(new_n696_), .C2(G36gat), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  INV_X1    g509(.A(G43gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n701_), .B2(new_n356_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT110), .Z(new_n713_));
  NAND4_X1  g512(.A1(new_n679_), .A2(G43gat), .A3(new_n685_), .A4(new_n355_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT47), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n714_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1330gat));
  INV_X1    g518(.A(G50gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n557_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n563_), .A2(new_n432_), .A3(new_n690_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n686_), .A2(new_n721_), .B1(new_n720_), .B2(new_n722_), .ZN(G1331gat));
  OAI21_X1  g522(.A(new_n301_), .B1(new_n621_), .B2(new_n561_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n270_), .A2(new_n614_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n552_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n270_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n724_), .B2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n655_), .A2(KEYINPUT111), .A3(new_n301_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n607_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n552_), .A2(G57gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n728_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT112), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n727_), .B2(new_n544_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n544_), .A2(G64gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n734_), .B2(new_n740_), .ZN(G1333gat));
  OR2_X1    g540(.A1(new_n356_), .A2(G71gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n725_), .A2(new_n355_), .A3(new_n726_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT49), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(G71gat), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n743_), .B2(G71gat), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n734_), .A2(new_n742_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750_));
  OAI221_X1 g549(.A(new_n750_), .B1(new_n746_), .B2(new_n747_), .C1(new_n734_), .C2(new_n742_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1334gat));
  OAI21_X1  g551(.A(G78gat), .B1(new_n727_), .B2(new_n557_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT50), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n432_), .A2(new_n203_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n734_), .B2(new_n755_), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n729_), .A2(new_n300_), .A3(new_n676_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n673_), .A2(KEYINPUT43), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n655_), .A2(new_n674_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n552_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n733_), .A2(new_n690_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n552_), .A2(G85gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n762_), .B2(new_n544_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n544_), .A2(G92gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n764_), .B2(new_n768_), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n762_), .B2(new_n356_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n356_), .A2(new_n245_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n731_), .A2(new_n690_), .A3(new_n732_), .A4(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT114), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(KEYINPUT114), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n770_), .B(new_n777_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1338gat));
  NOR2_X1   g578(.A1(new_n557_), .A2(G106gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n733_), .A2(new_n690_), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n220_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n761_), .B2(new_n432_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n781_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n784_), .A2(new_n786_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT53), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n784_), .A2(new_n786_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n784_), .A2(new_n786_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .A4(new_n781_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(G1339gat));
  NOR2_X1   g593(.A1(new_n300_), .A2(new_n606_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n268_), .A2(new_n269_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT116), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n268_), .A2(new_n798_), .A3(new_n795_), .A4(new_n269_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n589_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(new_n589_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n300_), .A2(new_n265_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n253_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n244_), .A2(new_n250_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n254_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n244_), .A2(new_n250_), .A3(KEYINPUT55), .A4(new_n252_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n806_), .B1(new_n253_), .B2(new_n807_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n262_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT56), .B(new_n262_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n805_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n294_), .A2(new_n297_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n293_), .A2(new_n286_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n297_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT118), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n266_), .A2(new_n819_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n689_), .B1(new_n818_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n823_), .A2(new_n265_), .A3(new_n819_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n817_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n253_), .A2(new_n807_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT117), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(new_n808_), .A3(new_n810_), .A4(new_n811_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n262_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n828_), .B1(new_n829_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT58), .B(new_n828_), .C1(new_n829_), .C2(new_n833_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n590_), .A3(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT57), .B(new_n689_), .C1(new_n818_), .C2(new_n824_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n827_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n804_), .B1(new_n840_), .B2(new_n606_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n841_), .A2(new_n552_), .A3(new_n560_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n300_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n606_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n804_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n550_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n849_), .B2(new_n560_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n842_), .A2(KEYINPUT59), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n301_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n844_), .B1(new_n852_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n729_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n842_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n729_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n854_), .ZN(G1341gat));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n842_), .A2(new_n859_), .A3(new_n676_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n606_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n859_), .ZN(G1342gat));
  INV_X1    g661(.A(G134gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n842_), .A2(new_n863_), .A3(new_n586_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n589_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1343gat));
  AOI21_X1  g665(.A(new_n552_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n557_), .A2(new_n355_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n544_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT119), .B1(new_n867_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n841_), .A2(new_n872_), .A3(new_n552_), .A4(new_n869_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n300_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G141gat), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n362_), .B(new_n300_), .C1(new_n871_), .C2(new_n873_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1344gat));
  OAI21_X1  g676(.A(new_n270_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G148gat), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n363_), .B(new_n270_), .C1(new_n871_), .C2(new_n873_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1345gat));
  OAI21_X1  g680(.A(new_n676_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n883_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n676_), .B(new_n885_), .C1(new_n871_), .C2(new_n873_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1346gat));
  INV_X1    g686(.A(G162gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n586_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n872_), .B1(new_n849_), .B2(new_n869_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n867_), .A2(KEYINPUT119), .A3(new_n870_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n672_), .A2(G162gat), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n888_), .A2(new_n889_), .B1(new_n892_), .B2(new_n893_), .ZN(G1347gat));
  NOR4_X1   g693(.A1(new_n841_), .A2(new_n550_), .A3(new_n544_), .A4(new_n558_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n300_), .A2(new_n315_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT120), .Z(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n550_), .A2(new_n544_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n848_), .A2(new_n300_), .A3(new_n559_), .A4(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n900_), .A2(new_n901_), .A3(G169gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n900_), .B2(G169gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n898_), .B1(new_n902_), .B2(new_n903_), .ZN(G1348gat));
  OR2_X1    g703(.A1(new_n317_), .A2(KEYINPUT121), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n317_), .A2(KEYINPUT121), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n895_), .A2(new_n270_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n895_), .A2(new_n270_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n906_), .ZN(G1349gat));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910_));
  INV_X1    g709(.A(new_n331_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n895_), .A2(new_n910_), .A3(new_n911_), .A4(new_n676_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n895_), .A2(new_n911_), .A3(new_n676_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT122), .ZN(new_n914_));
  AOI21_X1  g713(.A(G183gat), .B1(new_n895_), .B2(new_n676_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n912_), .B1(new_n914_), .B2(new_n915_), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n895_), .A2(new_n332_), .A3(new_n586_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n848_), .A2(new_n559_), .A3(new_n590_), .A4(new_n899_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n918_), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(KEYINPUT123), .B1(new_n918_), .B2(G190gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n917_), .B1(new_n919_), .B2(new_n920_), .ZN(G1351gat));
  NAND4_X1  g720(.A1(new_n848_), .A2(new_n300_), .A3(new_n868_), .A4(new_n899_), .ZN(new_n922_));
  INV_X1    g721(.A(G197gat), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n922_), .A2(KEYINPUT124), .A3(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n922_), .B2(new_n923_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n922_), .A2(new_n923_), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(G1352gat));
  AND3_X1   g726(.A1(new_n848_), .A2(new_n868_), .A3(new_n899_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n270_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g729(.A1(new_n848_), .A2(new_n676_), .A3(new_n868_), .A4(new_n899_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT63), .B(G211gat), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n934_));
  INV_X1    g733(.A(G211gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n931_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(KEYINPUT125), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n931_), .A2(new_n938_), .A3(new_n934_), .A4(new_n935_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n933_), .B1(new_n937_), .B2(new_n939_), .ZN(G1354gat));
  AND3_X1   g739(.A1(new_n928_), .A2(G218gat), .A3(new_n590_), .ZN(new_n941_));
  AND4_X1   g740(.A1(new_n586_), .A2(new_n848_), .A3(new_n868_), .A4(new_n899_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(G218gat), .B1(new_n942_), .B2(new_n943_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n941_), .B1(new_n944_), .B2(new_n945_), .ZN(G1355gat));
endmodule


