//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT12), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(G99gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(new_n205_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(KEYINPUT9), .A3(new_n212_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n206_), .A2(new_n211_), .A3(new_n213_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G85gat), .B(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT64), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n223_), .A2(new_n209_), .A3(new_n210_), .A4(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n216_), .A2(KEYINPUT65), .A3(new_n212_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n222_), .A2(new_n225_), .A3(new_n229_), .A4(new_n226_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n219_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT66), .B(G71gat), .ZN(new_n232_));
  INV_X1    g031(.A(G78gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n232_), .B(G78gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n203_), .B1(new_n231_), .B2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n231_), .A2(new_n241_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n228_), .A2(KEYINPUT67), .A3(new_n230_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n218_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT67), .B1(new_n228_), .B2(new_n230_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n241_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT12), .ZN(new_n249_));
  OAI221_X1 g048(.A(new_n202_), .B1(new_n242_), .B2(new_n243_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT68), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n247_), .A2(new_n249_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n242_), .A2(new_n243_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .A4(new_n202_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n231_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(new_n248_), .ZN(new_n257_));
  OAI211_X1 g056(.A(G230gat), .B(G233gat), .C1(new_n257_), .C2(new_n243_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n255_), .A3(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G120gat), .B(G148gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G176gat), .B(G204gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n262_), .B(new_n263_), .Z(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n251_), .A2(new_n255_), .A3(new_n258_), .A4(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT13), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT13), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT73), .B(G8gat), .Z(new_n273_));
  INV_X1    g072(.A(G1gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT14), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G15gat), .B(G22gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G1gat), .B(G8gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G29gat), .B(G36gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G43gat), .B(G50gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT15), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n282_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n284_), .B1(new_n279_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G229gat), .A2(G233gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n279_), .B(new_n285_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G113gat), .B(G141gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT74), .ZN(new_n292_));
  XOR2_X1   g091(.A(G169gat), .B(G197gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n290_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n272_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n299_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n303_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312_));
  INV_X1    g111(.A(G169gat), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT24), .B1(new_n315_), .B2(new_n300_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT78), .B1(new_n316_), .B2(new_n308_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT25), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(KEYINPUT75), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT76), .B(G190gat), .Z(new_n326_));
  OAI211_X1 g125(.A(new_n319_), .B(new_n325_), .C1(new_n326_), .C2(new_n318_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n315_), .A2(KEYINPUT24), .A3(new_n328_), .A4(new_n300_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n311_), .A2(new_n317_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT21), .ZN(new_n331_));
  INV_X1    g130(.A(G197gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(G204gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(G204gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n331_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G218gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G211gat), .ZN(new_n340_));
  INV_X1    g139(.A(G211gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G218gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n342_), .A3(KEYINPUT88), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n335_), .A2(new_n334_), .ZN(new_n348_));
  INV_X1    g147(.A(G204gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G197gat), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n348_), .A2(new_n331_), .A3(new_n337_), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n335_), .A2(new_n350_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n343_), .B1(KEYINPUT21), .B2(new_n352_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n338_), .A2(new_n347_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n328_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G169gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n356_), .B2(new_n314_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n326_), .A2(G183gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(new_n308_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n330_), .A2(new_n354_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT26), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n320_), .A2(G183gat), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n319_), .A2(new_n362_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n315_), .A2(new_n328_), .A3(new_n300_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n315_), .A2(new_n300_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n308_), .B1(new_n369_), .B2(new_n367_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(KEYINPUT90), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT90), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n369_), .A2(new_n367_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(new_n308_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n309_), .B1(G183gat), .B2(G190gat), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n371_), .A2(new_n374_), .B1(new_n357_), .B2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT20), .B(new_n360_), .C1(new_n376_), .C2(new_n354_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT19), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n377_), .A2(KEYINPUT97), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT97), .B1(new_n377_), .B2(new_n379_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n354_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n330_), .A2(new_n359_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n354_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n383_), .A2(KEYINPUT20), .A3(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n380_), .B(new_n381_), .C1(new_n382_), .C2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT18), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(KEYINPUT32), .A3(new_n392_), .ZN(new_n393_));
  OAI22_X1  g192(.A1(KEYINPUT83), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT2), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT2), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(G141gat), .A3(G148gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT83), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n396_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT84), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n396_), .A2(new_n401_), .A3(new_n405_), .A4(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G155gat), .A2(G162gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G127gat), .B(G134gat), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT80), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G127gat), .B(G134gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G113gat), .B(G120gat), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n415_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(G141gat), .A2(G148gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n397_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n408_), .B1(new_n410_), .B2(KEYINPUT1), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT82), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n408_), .A2(KEYINPUT1), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(KEYINPUT82), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n425_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n413_), .A2(new_n423_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n415_), .A2(new_n418_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n419_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n415_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n411_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(new_n432_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n434_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n434_), .A2(new_n440_), .A3(KEYINPUT4), .ZN(new_n443_));
  INV_X1    g242(.A(new_n441_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n440_), .B2(KEYINPUT4), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n442_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT0), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G57gat), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n447_), .A2(KEYINPUT0), .ZN(new_n450_));
  INV_X1    g249(.A(G57gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(KEYINPUT0), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n449_), .A2(new_n453_), .A3(G85gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(G85gat), .B1(new_n449_), .B2(new_n453_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n446_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n442_), .B(new_n458_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n377_), .A2(new_n379_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT91), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT91), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n377_), .A2(new_n463_), .A3(new_n379_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n383_), .A2(KEYINPUT20), .A3(new_n382_), .A4(new_n386_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n393_), .A2(new_n460_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n434_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n456_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n470_), .B2(new_n456_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n441_), .B1(new_n440_), .B2(KEYINPUT4), .ZN(new_n474_));
  OAI22_X1  g273(.A1(new_n472_), .A2(new_n473_), .B1(new_n443_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT96), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n459_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n459_), .B2(new_n478_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  OAI22_X1  g280(.A1(new_n479_), .A2(new_n480_), .B1(new_n481_), .B2(new_n459_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n392_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n377_), .A2(new_n463_), .A3(new_n379_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n463_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n392_), .B(new_n466_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n484_), .B1(new_n485_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n466_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n392_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(KEYINPUT92), .A3(new_n488_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n469_), .B1(new_n483_), .B2(new_n495_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n439_), .A2(KEYINPUT29), .A3(new_n432_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(KEYINPUT85), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT28), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n439_), .A2(new_n432_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT29), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(KEYINPUT85), .A3(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n503_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT28), .B1(new_n505_), .B2(new_n498_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G78gat), .B(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT29), .B1(new_n439_), .B2(new_n432_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G228gat), .A2(G233gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n354_), .B2(KEYINPUT86), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n510_), .A2(new_n385_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n510_), .B2(new_n385_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n509_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n385_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n512_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n510_), .A2(new_n512_), .A3(new_n385_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n508_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G22gat), .B(G50gat), .Z(new_n521_));
  AND3_X1   g320(.A1(new_n515_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n515_), .B2(new_n520_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n507_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n521_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n513_), .A2(new_n514_), .A3(new_n509_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n508_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n504_), .A2(new_n506_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n515_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G71gat), .B(G99gat), .ZN(new_n535_));
  INV_X1    g334(.A(G43gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G227gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(G15gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n537_), .B(new_n540_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n330_), .A2(KEYINPUT30), .A3(new_n359_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT30), .B1(new_n330_), .B2(new_n359_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n384_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n537_), .B(new_n540_), .Z(new_n547_));
  NAND3_X1  g346(.A1(new_n330_), .A2(KEYINPUT30), .A3(new_n359_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT81), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n544_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n438_), .B(KEYINPUT31), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT79), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n551_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n553_), .A2(new_n554_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n542_), .A2(new_n543_), .A3(new_n541_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n547_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT81), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n544_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n534_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n460_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n524_), .A2(new_n563_), .A3(new_n532_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n563_), .B1(new_n524_), .B2(new_n532_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n485_), .A2(new_n489_), .A3(KEYINPUT27), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n388_), .A2(new_n492_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n465_), .A2(KEYINPUT98), .A3(new_n392_), .A4(new_n466_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n488_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n570_), .B1(new_n575_), .B2(KEYINPUT27), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n496_), .A2(new_n565_), .B1(new_n569_), .B2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n298_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n283_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT70), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT70), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n587_), .B(new_n283_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT35), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n231_), .A2(new_n282_), .B1(new_n590_), .B2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n256_), .A2(new_n285_), .ZN(new_n595_));
  OAI211_X1 g394(.A(KEYINPUT35), .B(new_n592_), .C1(new_n595_), .C2(KEYINPUT71), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n589_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n584_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n582_), .A2(new_n583_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  OAI221_X1 g403(.A(new_n600_), .B1(new_n604_), .B2(new_n584_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n579_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n579_), .A3(new_n605_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n241_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n279_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(G127gat), .B(G155gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT17), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n613_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n613_), .A2(new_n619_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n609_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n578_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n274_), .A3(new_n460_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT99), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(KEYINPUT38), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n298_), .A2(new_n623_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n603_), .A2(new_n605_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n577_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n566_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n628_), .A2(KEYINPUT38), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT100), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT100), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n629_), .B(new_n636_), .C1(new_n638_), .C2(new_n639_), .ZN(G1324gat));
  INV_X1    g439(.A(new_n576_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G8gat), .B1(new_n635_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT39), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n626_), .A2(new_n273_), .A3(new_n576_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g445(.A(G15gat), .B1(new_n635_), .B2(new_n564_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT41), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n626_), .A2(new_n539_), .A3(new_n563_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(G1326gat));
  OAI21_X1  g450(.A(G22gat), .B1(new_n635_), .B2(new_n534_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT42), .ZN(new_n653_));
  INV_X1    g452(.A(G22gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n534_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n626_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n633_), .A2(new_n623_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n578_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n460_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n577_), .A2(new_n609_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n577_), .B2(new_n609_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n577_), .A2(new_n609_), .A3(KEYINPUT101), .A4(new_n662_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n624_), .A4(new_n298_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n669_), .A2(G29gat), .A3(new_n460_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n666_), .A2(new_n667_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n298_), .A2(new_n624_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n671_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n661_), .B1(new_n670_), .B2(new_n674_), .ZN(G1328gat));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n576_), .A3(new_n669_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n659_), .A2(G36gat), .A3(new_n641_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT45), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1329gat));
  NAND4_X1  g481(.A1(new_n674_), .A2(G43gat), .A3(new_n563_), .A4(new_n669_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n536_), .B1(new_n659_), .B2(new_n564_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT102), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g486(.A1(new_n674_), .A2(new_n655_), .A3(new_n669_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G50gat), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT103), .ZN(new_n690_));
  OR3_X1    g489(.A1(new_n659_), .A2(G50gat), .A3(new_n534_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1331gat));
  INV_X1    g491(.A(new_n272_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(new_n624_), .A3(new_n296_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n634_), .A2(new_n694_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n695_), .A2(new_n451_), .A3(new_n566_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT104), .Z(new_n697_));
  NOR2_X1   g496(.A1(new_n693_), .A2(new_n296_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n577_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n625_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n460_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n697_), .A2(new_n702_), .ZN(G1332gat));
  OAI21_X1  g502(.A(G64gat), .B1(new_n695_), .B2(new_n641_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT106), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT105), .B(KEYINPUT48), .Z(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n700_), .A2(G64gat), .A3(new_n641_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(G1333gat));
  OAI21_X1  g509(.A(G71gat), .B1(new_n695_), .B2(new_n564_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT49), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n564_), .A2(G71gat), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT107), .Z(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n700_), .B2(new_n714_), .ZN(G1334gat));
  OAI21_X1  g514(.A(G78gat), .B1(new_n695_), .B2(new_n534_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT50), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n701_), .A2(new_n233_), .A3(new_n655_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1335gat));
  NAND2_X1  g518(.A1(new_n698_), .A2(new_n624_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n566_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n699_), .A2(new_n658_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n214_), .A3(new_n460_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1336gat));
  AOI21_X1  g525(.A(G92gat), .B1(new_n724_), .B2(new_n576_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT108), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n641_), .A2(new_n215_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n721_), .B2(new_n729_), .ZN(G1337gat));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(KEYINPUT110), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n564_), .B(new_n720_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(new_n208_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n720_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n668_), .A2(new_n563_), .A3(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(KEYINPUT109), .A3(G99gat), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n563_), .A2(new_n204_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n724_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n734_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n743_), .ZN(new_n745_));
  AOI211_X1 g544(.A(KEYINPUT111), .B(new_n745_), .C1(new_n737_), .C2(new_n740_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n733_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n736_), .A2(new_n735_), .A3(new_n208_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT109), .B1(new_n739_), .B2(G99gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n743_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n741_), .A2(new_n734_), .A3(new_n743_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n732_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n747_), .A2(new_n753_), .ZN(G1338gat));
  AOI21_X1  g553(.A(new_n205_), .B1(new_n721_), .B2(new_n655_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n757_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n724_), .A2(new_n205_), .A3(new_n655_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g561(.A1(new_n607_), .A2(new_n608_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n272_), .A2(new_n296_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n623_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT113), .B1(new_n765_), .B2(KEYINPUT54), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n625_), .A2(new_n767_), .A3(new_n768_), .A4(new_n764_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(KEYINPUT54), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n766_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n250_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n202_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n251_), .A2(new_n255_), .A3(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n264_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n780_), .B(new_n266_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n294_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n267_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT115), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT58), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n782_), .A2(new_n787_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n763_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n296_), .A2(new_n267_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n268_), .A2(new_n785_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n632_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT119), .B1(new_n792_), .B2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n782_), .A2(new_n787_), .A3(new_n790_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n790_), .B1(new_n782_), .B2(new_n787_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n609_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n801_), .B(new_n802_), .C1(KEYINPUT57), .C2(new_n796_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n798_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n772_), .B1(new_n805_), .B2(new_n624_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n641_), .A2(new_n460_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n807_), .A2(new_n564_), .A3(new_n655_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT116), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n794_), .A2(new_n795_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT114), .B(new_n813_), .C1(new_n814_), .C2(new_n632_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n796_), .B2(KEYINPUT57), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n801_), .A2(new_n815_), .A3(new_n817_), .A4(new_n804_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n624_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n809_), .B1(new_n819_), .B2(new_n771_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  OAI22_X1  g620(.A1(new_n806_), .A2(new_n812_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822_), .B2(new_n297_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n820_), .B(KEYINPUT117), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n297_), .A2(G113gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n823_), .B1(new_n825_), .B2(new_n826_), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n822_), .B2(new_n693_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT60), .ZN(new_n829_));
  INV_X1    g628(.A(G120gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n272_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT120), .B1(new_n824_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n819_), .A2(new_n771_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n810_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n820_), .A2(new_n837_), .ZN(new_n838_));
  AND4_X1   g637(.A1(KEYINPUT120), .A2(new_n836_), .A3(new_n838_), .A4(new_n832_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n828_), .B1(new_n833_), .B2(new_n839_), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n822_), .B2(new_n624_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n624_), .A2(G127gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n825_), .B2(new_n842_), .ZN(G1342gat));
  AOI21_X1  g642(.A(G134gat), .B1(new_n824_), .B2(new_n632_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT121), .B(G134gat), .Z(new_n845_));
  NOR3_X1   g644(.A1(new_n822_), .A2(new_n763_), .A3(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1343gat));
  NAND2_X1  g646(.A1(new_n834_), .A2(new_n568_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n807_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n296_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n272_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT122), .B(G148gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  NAND2_X1  g653(.A1(new_n849_), .A2(new_n623_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  INV_X1    g656(.A(G162gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n849_), .A2(new_n858_), .A3(new_n632_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n848_), .A2(new_n763_), .A3(new_n807_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n858_), .B2(new_n860_), .ZN(G1347gat));
  NAND2_X1  g660(.A1(new_n576_), .A2(new_n566_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n563_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT123), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n655_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n806_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(new_n296_), .A3(new_n356_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n792_), .A2(new_n797_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n870_), .A2(new_n802_), .B1(KEYINPUT57), .B2(new_n796_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n623_), .B1(new_n871_), .B2(new_n798_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n296_), .B(new_n866_), .C1(new_n872_), .C2(new_n772_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n873_), .A2(new_n874_), .A3(G169gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(G169gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n869_), .B1(new_n875_), .B2(new_n876_), .ZN(G1348gat));
  NOR3_X1   g676(.A1(new_n806_), .A2(new_n693_), .A3(new_n867_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT124), .B1(new_n878_), .B2(G176gat), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n272_), .B(new_n866_), .C1(new_n872_), .C2(new_n772_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n881_), .A3(new_n314_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n655_), .B1(new_n819_), .B2(new_n771_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n865_), .A2(new_n314_), .A3(new_n693_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n879_), .A2(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1349gat));
  AOI21_X1  g684(.A(new_n624_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n866_), .B(new_n886_), .C1(new_n872_), .C2(new_n772_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n865_), .A2(new_n624_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n883_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(G183gat), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n887_), .B(KEYINPUT125), .C1(G183gat), .C2(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1350gat));
  NAND4_X1  g693(.A1(new_n868_), .A2(new_n632_), .A3(new_n319_), .A4(new_n362_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n806_), .A2(new_n763_), .A3(new_n867_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n361_), .ZN(G1351gat));
  NAND4_X1  g696(.A1(new_n834_), .A2(new_n296_), .A3(new_n568_), .A4(new_n863_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(new_n899_), .A3(new_n332_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n332_), .B2(new_n898_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n898_), .B2(new_n332_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1352gat));
  NOR2_X1   g702(.A1(new_n848_), .A2(new_n862_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n272_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g705(.A1(new_n834_), .A2(new_n568_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT63), .B(G211gat), .Z(new_n908_));
  NAND4_X1  g707(.A1(new_n907_), .A2(new_n623_), .A3(new_n863_), .A4(new_n908_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n834_), .A2(new_n623_), .A3(new_n568_), .A4(new_n863_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(new_n341_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n909_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1354gat));
  NAND3_X1  g715(.A1(new_n904_), .A2(new_n339_), .A3(new_n632_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n848_), .A2(new_n763_), .A3(new_n862_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n339_), .B2(new_n918_), .ZN(G1355gat));
endmodule


