//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT85), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT85), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n207_), .A2(new_n204_), .A3(G183gat), .A4(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT84), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(G183gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n206_), .A2(new_n208_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT86), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT86), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n206_), .A2(new_n214_), .A3(new_n217_), .A4(new_n208_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT26), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G190gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G169gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n222_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n203_), .A2(new_n205_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n229_), .A2(new_n232_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n224_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT30), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n239_), .A2(KEYINPUT88), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT87), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G15gat), .B(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n240_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT91), .ZN(new_n248_));
  INV_X1    g047(.A(G134gat), .ZN(new_n249_));
  INV_X1    g048(.A(G120gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G113gat), .ZN(new_n251_));
  INV_X1    g050(.A(G113gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G120gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n255_), .A2(new_n256_), .A3(G127gat), .ZN(new_n257_));
  INV_X1    g056(.A(G127gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n252_), .A2(G120gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n250_), .A2(G113gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT90), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n249_), .B1(new_n257_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(G127gat), .B1(new_n255_), .B2(new_n256_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n258_), .A3(new_n262_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(G134gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT31), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n248_), .B1(new_n270_), .B2(KEYINPUT89), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n239_), .A2(KEYINPUT88), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n246_), .B1(new_n240_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n247_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n248_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n247_), .A2(new_n275_), .A3(new_n273_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n276_), .B2(new_n271_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT0), .ZN(new_n280_));
  INV_X1    g079(.A(G57gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(G85gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(G155gat), .A3(G162gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT93), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n284_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n285_), .A2(KEYINPUT93), .A3(G155gat), .A4(G162gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT92), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(KEYINPUT1), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n291_), .A2(new_n290_), .A3(KEYINPUT1), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n288_), .B(new_n289_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G141gat), .B(G148gat), .Z(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n284_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n291_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT3), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(G141gat), .B2(G148gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n298_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n296_), .A2(new_n308_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n265_), .A2(G134gat), .A3(new_n266_), .ZN(new_n310_));
  AOI21_X1  g109(.A(G134gat), .B1(new_n265_), .B2(new_n266_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT99), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n307_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n264_), .A2(new_n267_), .A3(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n268_), .A2(KEYINPUT99), .A3(new_n309_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT4), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT100), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n312_), .B2(KEYINPUT4), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n314_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT100), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n318_), .A2(new_n320_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n283_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n320_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n312_), .A2(new_n321_), .A3(KEYINPUT4), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT100), .B1(new_n323_), .B2(new_n324_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n324_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n328_), .B(new_n283_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n329_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G218gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G211gat), .ZN(new_n342_));
  INV_X1    g141(.A(G211gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G218gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT21), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n342_), .A2(new_n344_), .A3(KEYINPUT21), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n348_), .A2(KEYINPUT21), .A3(new_n342_), .A4(new_n344_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n314_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(G228gat), .A3(G233gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n353_), .B(new_n357_), .C1(new_n314_), .C2(new_n354_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n340_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n358_), .A3(new_n340_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n314_), .A2(new_n354_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G22gat), .B(G50gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n363_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT95), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n359_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n360_), .A2(new_n368_), .A3(new_n361_), .A4(new_n367_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT18), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G64gat), .ZN(new_n375_));
  INV_X1    g174(.A(G92gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n238_), .A2(new_n353_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n230_), .A2(KEYINPUT22), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G169gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n382_), .A3(new_n222_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n219_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n203_), .A2(new_n205_), .B1(new_n213_), .B2(new_n209_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n234_), .A2(KEYINPUT96), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT96), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT24), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n389_), .A3(new_n233_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n231_), .A2(new_n219_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n213_), .A2(KEYINPUT25), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT25), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G183gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n209_), .A2(KEYINPUT26), .ZN(new_n397_));
  AND4_X1   g196(.A1(new_n227_), .A2(new_n394_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n206_), .A2(new_n208_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n386_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n351_), .A2(new_n352_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n379_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT97), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT19), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n378_), .A2(new_n404_), .A3(new_n405_), .A4(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n213_), .A2(new_n209_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n236_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n223_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n388_), .A2(KEYINPUT24), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n234_), .A2(KEYINPUT96), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n231_), .B(new_n219_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT26), .B(G190gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n228_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n417_), .A3(new_n390_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n412_), .B1(new_n418_), .B2(new_n400_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n379_), .B1(new_n419_), .B2(new_n353_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n224_), .A2(new_n403_), .A3(new_n237_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n407_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT20), .B(new_n408_), .C1(new_n419_), .C2(new_n353_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n403_), .B1(new_n224_), .B2(new_n237_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT97), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n377_), .A2(new_n409_), .A3(new_n423_), .A4(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n375_), .B(G92gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT102), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n422_), .A2(new_n407_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n408_), .B1(new_n378_), .B2(new_n404_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT27), .B(new_n427_), .C1(new_n429_), .C2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n409_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n428_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n427_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NOR4_X1   g238(.A1(new_n278_), .A2(new_n338_), .A3(new_n372_), .A4(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n335_), .A2(KEYINPUT33), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n327_), .A2(new_n442_), .A3(new_n328_), .A4(new_n283_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n330_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n319_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n283_), .B1(new_n318_), .B2(new_n330_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n436_), .A2(KEYINPUT98), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT98), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n435_), .A2(new_n449_), .A3(new_n427_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n444_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n377_), .A2(KEYINPUT32), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT101), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n452_), .B(new_n432_), .C1(new_n453_), .C2(new_n434_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n434_), .A2(KEYINPUT101), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n329_), .B2(new_n336_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n372_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n337_), .A2(new_n372_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(new_n439_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n278_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT103), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT103), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n463_), .B(new_n278_), .C1(new_n458_), .C2(new_n460_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n440_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT79), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G229gat), .A2(G233gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G29gat), .B(G36gat), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n470_), .A2(KEYINPUT69), .ZN(new_n471_));
  INV_X1    g270(.A(G43gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(KEYINPUT69), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G50gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G8gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT72), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT71), .B(G1gat), .Z(new_n482_));
  INV_X1    g281(.A(G8gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT14), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n480_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n470_), .B(KEYINPUT69), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G43gat), .ZN(new_n491_));
  AOI21_X1  g290(.A(G50gat), .B1(new_n491_), .B2(new_n474_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n478_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n476_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(G50gat), .A3(new_n474_), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n494_), .A2(new_n495_), .B1(new_n488_), .B2(new_n487_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n469_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT77), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT77), .B(new_n469_), .C1(new_n493_), .C2(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(new_n478_), .B2(new_n492_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n494_), .A2(KEYINPUT15), .A3(new_n495_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n493_), .B1(new_n505_), .B2(new_n489_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT78), .B1(new_n506_), .B2(new_n468_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n489_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n510_));
  NOR4_X1   g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n493_), .A4(new_n469_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n467_), .B(new_n501_), .C1(new_n507_), .C2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G169gat), .B(G197gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G141gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT80), .B(G113gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT81), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n478_), .A2(new_n492_), .A3(new_n502_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT15), .B1(new_n494_), .B2(new_n495_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n489_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n493_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n468_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n510_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n506_), .A2(KEYINPUT78), .A3(new_n468_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n467_), .B1(new_n526_), .B2(new_n501_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n466_), .B1(new_n518_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n501_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT79), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n530_), .A2(KEYINPUT82), .A3(new_n517_), .A4(new_n512_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n526_), .A2(new_n501_), .A3(new_n516_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT83), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT83), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n528_), .A2(new_n531_), .A3(new_n535_), .A4(new_n532_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n465_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT6), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n541_));
  OR3_X1    g340(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G85gat), .B(G92gat), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT8), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT66), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n540_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n544_), .B2(new_n552_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT65), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT10), .B(G99gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(G106gat), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n556_), .A2(KEYINPUT65), .A3(G106gat), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n550_), .B(new_n554_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n543_), .A2(KEYINPUT8), .A3(new_n544_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n547_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n505_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n494_), .A2(new_n495_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  OAI22_X1  g366(.A1(new_n565_), .A2(new_n563_), .B1(KEYINPUT35), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n567_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT35), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n564_), .B(new_n569_), .C1(new_n572_), .C2(new_n571_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n577_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n574_), .A2(new_n576_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(KEYINPUT36), .A3(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(KEYINPUT37), .A3(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G57gat), .B(G64gat), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n591_), .A2(KEYINPUT11), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(KEYINPUT11), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G71gat), .B(G78gat), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(new_n594_), .A3(KEYINPUT11), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n563_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n596_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n599_), .A2(new_n547_), .A3(new_n561_), .A4(new_n562_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(KEYINPUT12), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n563_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT64), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n598_), .A2(new_n600_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT68), .ZN(new_n613_));
  XOR2_X1   g412(.A(G120gat), .B(G148gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n615_), .B(new_n616_), .Z(new_n617_));
  NAND2_X1  g416(.A1(new_n611_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n608_), .A2(new_n610_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT13), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT73), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n599_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n489_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT17), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(KEYINPUT17), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n634_), .B(KEYINPUT76), .Z(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n628_), .B2(KEYINPUT74), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT74), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n627_), .A2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n623_), .A2(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n538_), .A2(new_n590_), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n338_), .A3(new_n482_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT38), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n465_), .A2(new_n586_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n533_), .A2(KEYINPUT104), .A3(new_n622_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT104), .B1(new_n533_), .B2(new_n622_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(new_n641_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT105), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n337_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n645_), .A2(new_n652_), .ZN(G1324gat));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n646_), .A2(new_n439_), .A3(new_n649_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(G8gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G8gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n661_));
  INV_X1    g460(.A(new_n439_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(G8gat), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n660_), .A2(new_n661_), .B1(new_n643_), .B2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(KEYINPUT107), .A2(KEYINPUT39), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n655_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n656_), .A2(G8gat), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT106), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n656_), .A2(new_n657_), .A3(G8gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n661_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n643_), .A2(new_n663_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(KEYINPUT108), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n654_), .B1(new_n667_), .B2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n664_), .A2(new_n655_), .A3(new_n666_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(KEYINPUT108), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(KEYINPUT40), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(G1325gat));
  INV_X1    g478(.A(new_n643_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n680_), .A2(G15gat), .A3(new_n278_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n651_), .A2(new_n278_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT41), .B1(new_n682_), .B2(G15gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(new_n372_), .ZN(new_n686_));
  OR3_X1    g485(.A1(new_n680_), .A2(G22gat), .A3(new_n686_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n651_), .A2(new_n686_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(new_n689_), .A3(G22gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G22gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1327gat));
  NAND3_X1  g491(.A1(new_n586_), .A2(new_n622_), .A3(new_n641_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n465_), .A2(new_n537_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n338_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n641_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n647_), .A2(new_n648_), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n465_), .B2(new_n590_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n465_), .A2(KEYINPUT43), .A3(new_n590_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(KEYINPUT109), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n465_), .A2(new_n701_), .A3(KEYINPUT43), .A4(new_n590_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n697_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n703_), .A2(G29gat), .A3(new_n338_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n462_), .A2(new_n464_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n440_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  INV_X1    g507(.A(new_n590_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n701_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n699_), .A2(KEYINPUT109), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n698_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT44), .B1(new_n713_), .B2(new_n697_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n695_), .B1(new_n704_), .B2(new_n715_), .ZN(G1328gat));
  NAND2_X1  g515(.A1(new_n703_), .A2(new_n439_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G36gat), .B1(new_n717_), .B2(new_n714_), .ZN(new_n718_));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n694_), .A2(new_n719_), .A3(new_n439_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT45), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT46), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT110), .B(new_n725_), .C1(new_n718_), .C2(new_n721_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1329gat));
  NAND3_X1  g526(.A1(new_n703_), .A2(G43gat), .A3(new_n277_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n694_), .A2(new_n277_), .ZN(new_n729_));
  OAI22_X1  g528(.A1(new_n728_), .A2(new_n714_), .B1(G43gat), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g530(.A(G50gat), .B1(new_n694_), .B2(new_n372_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n703_), .A2(G50gat), .A3(new_n372_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n715_), .ZN(G1331gat));
  NOR2_X1   g533(.A1(new_n622_), .A2(new_n641_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n646_), .A2(new_n537_), .A3(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n337_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n533_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n590_), .A2(new_n738_), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n707_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n338_), .A2(new_n281_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n736_), .B2(new_n662_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n662_), .A2(G64gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n740_), .B2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n736_), .B2(new_n278_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n278_), .A2(G71gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n740_), .B2(new_n750_), .ZN(G1334gat));
  OAI21_X1  g550(.A(G78gat), .B1(new_n736_), .B2(new_n686_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT50), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n686_), .A2(G78gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n740_), .B2(new_n754_), .ZN(G1335gat));
  NAND3_X1  g554(.A1(new_n738_), .A2(new_n641_), .A3(new_n623_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n585_), .B2(new_n583_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n707_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(G85gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n338_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n756_), .B(KEYINPUT112), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n713_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n713_), .A2(KEYINPUT113), .A3(new_n763_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n337_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n761_), .B1(new_n768_), .B2(new_n760_), .ZN(G1336gat));
  OAI21_X1  g568(.A(new_n376_), .B1(new_n758_), .B2(new_n662_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT114), .Z(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(new_n767_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n439_), .A2(G92gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT115), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n772_), .B2(new_n774_), .ZN(G1337gat));
  NAND3_X1  g574(.A1(new_n759_), .A2(new_n557_), .A3(new_n277_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n278_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n777_));
  INV_X1    g576(.A(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT51), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n776_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1338gat));
  OAI211_X1 g582(.A(new_n372_), .B(new_n763_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT117), .B1(new_n784_), .B2(G106gat), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n784_), .A2(KEYINPUT117), .A3(G106gat), .ZN(new_n787_));
  XOR2_X1   g586(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n787_), .A2(new_n789_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n759_), .A2(new_n558_), .A3(new_n372_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n789_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n785_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n793_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n794_), .A2(new_n798_), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n439_), .A2(new_n337_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n278_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n604_), .A2(new_n607_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n608_), .A2(KEYINPUT55), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n604_), .A2(new_n806_), .A3(new_n607_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n803_), .B(KEYINPUT56), .C1(new_n808_), .C2(new_n619_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n620_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n806_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT55), .B(new_n606_), .C1(new_n601_), .C2(new_n603_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n617_), .B1(new_n813_), .B2(new_n804_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n814_), .B2(new_n803_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n810_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n533_), .A2(new_n816_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n493_), .A2(new_n496_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n516_), .B1(new_n818_), .B2(new_n468_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n506_), .A2(new_n469_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n532_), .A2(new_n621_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n586_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT57), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT121), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n826_), .A3(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n532_), .A2(new_n620_), .A3(new_n821_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT119), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n532_), .A2(new_n831_), .A3(new_n620_), .A4(new_n821_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n814_), .B(KEYINPUT56), .Z(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(KEYINPUT120), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(KEYINPUT120), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n834_), .A3(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n709_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841_));
  INV_X1    g640(.A(new_n822_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n533_), .B2(new_n816_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(new_n586_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n840_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n696_), .B1(new_n828_), .B2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n590_), .A2(new_n536_), .A3(new_n534_), .A4(new_n642_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n686_), .B(new_n802_), .C1(new_n846_), .C2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n252_), .A3(new_n533_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n826_), .B1(new_n823_), .B2(KEYINPUT57), .ZN(new_n855_));
  NOR4_X1   g654(.A1(new_n843_), .A2(KEYINPUT121), .A3(new_n841_), .A4(new_n586_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n844_), .B(new_n840_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n641_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n849_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n372_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n854_), .B1(new_n860_), .B2(new_n802_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n849_), .B1(new_n857_), .B2(new_n641_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n802_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n862_), .A2(KEYINPUT59), .A3(new_n372_), .A4(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n853_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n860_), .A2(new_n854_), .A3(new_n802_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(KEYINPUT122), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n537_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n852_), .B1(new_n869_), .B2(new_n252_), .ZN(G1340gat));
  NAND3_X1  g669(.A1(new_n866_), .A2(new_n623_), .A3(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT123), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n866_), .A2(new_n867_), .A3(new_n873_), .A4(new_n623_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(G120gat), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n622_), .B2(G120gat), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n851_), .B(new_n877_), .C1(new_n876_), .C2(G120gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(G1341gat));
  NAND3_X1  g678(.A1(new_n851_), .A2(new_n258_), .A3(new_n696_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n641_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n258_), .ZN(G1342gat));
  NAND3_X1  g681(.A1(new_n851_), .A2(new_n249_), .A3(new_n586_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n590_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n249_), .ZN(G1343gat));
  NOR4_X1   g684(.A1(new_n862_), .A2(new_n686_), .A3(new_n277_), .A4(new_n801_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n533_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT124), .B(G141gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1344gat));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n623_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g690(.A1(new_n886_), .A2(new_n696_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  INV_X1    g693(.A(G162gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n886_), .A2(new_n895_), .A3(new_n586_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n886_), .A2(new_n709_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(G1347gat));
  NAND2_X1  g697(.A1(new_n858_), .A2(new_n859_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n686_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n277_), .A2(new_n337_), .A3(new_n439_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G169gat), .B1(new_n902_), .B2(new_n738_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT62), .B(G169gat), .C1(new_n902_), .C2(new_n738_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n900_), .A2(new_n901_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(new_n221_), .A3(new_n533_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n905_), .A2(new_n906_), .A3(new_n908_), .ZN(G1348gat));
  AND2_X1   g708(.A1(new_n222_), .A2(KEYINPUT125), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT125), .B(G176gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n907_), .A2(new_n623_), .ZN(new_n912_));
  MUX2_X1   g711(.A(new_n910_), .B(new_n911_), .S(new_n912_), .Z(G1349gat));
  NAND2_X1  g712(.A1(new_n907_), .A2(new_n696_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n228_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n213_), .B2(new_n914_), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n902_), .B2(new_n590_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n907_), .A2(new_n586_), .A3(new_n416_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1351gat));
  NOR4_X1   g718(.A1(new_n862_), .A2(new_n459_), .A3(new_n662_), .A4(new_n277_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n533_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT126), .B(G197gat), .Z(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1352gat));
  NAND2_X1  g722(.A1(new_n920_), .A2(new_n623_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g724(.A1(new_n920_), .A2(new_n696_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  AND2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n926_), .B2(new_n927_), .ZN(G1354gat));
  AOI21_X1  g729(.A(G218gat), .B1(new_n920_), .B2(new_n586_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n709_), .A2(G218gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT127), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n920_), .B2(new_n933_), .ZN(G1355gat));
endmodule


