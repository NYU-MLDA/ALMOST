//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT68), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n215_), .A2(new_n217_), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT65), .B(KEYINPUT8), .Z(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT10), .B(G99gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n212_), .A2(new_n213_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT64), .B(G92gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(G85gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .A4(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G29gat), .B(G36gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G43gat), .B(G50gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n233_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n231_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  OAI221_X1 g036(.A(new_n205_), .B1(KEYINPUT35), .B2(new_n203_), .C1(new_n230_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n218_), .B(KEYINPUT66), .C1(new_n219_), .C2(new_n220_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n220_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n244_), .A3(new_n229_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT67), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n240_), .A2(new_n244_), .A3(new_n247_), .A4(new_n229_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n237_), .B(KEYINPUT15), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n204_), .B(new_n239_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n252_));
  OAI211_X1 g051(.A(KEYINPUT35), .B(new_n203_), .C1(new_n252_), .C2(new_n238_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G190gat), .B(G218gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G134gat), .B(G162gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT36), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n251_), .A2(new_n253_), .A3(KEYINPUT69), .A4(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n251_), .A2(new_n253_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n256_), .B(KEYINPUT36), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT37), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n269_), .A3(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G127gat), .B(G155gat), .ZN(new_n273_));
  INV_X1    g072(.A(G211gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT16), .B(G183gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G1gat), .A2(G8gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT14), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G1gat), .B(G8gat), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT70), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n285_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G57gat), .B(G64gat), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(KEYINPUT11), .ZN(new_n291_));
  XOR2_X1   g090(.A(G71gat), .B(G78gat), .Z(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n291_), .A2(new_n292_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n288_), .B(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n277_), .B1(new_n297_), .B2(KEYINPUT17), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(KEYINPUT17), .B2(new_n277_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n297_), .A2(KEYINPUT71), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n272_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(KEYINPUT12), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G230gat), .A2(G233gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n221_), .A2(new_n295_), .A3(new_n229_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n295_), .B1(new_n229_), .B2(new_n221_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(KEYINPUT12), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n305_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n309_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n306_), .B1(new_n312_), .B2(new_n308_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G120gat), .B(G148gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(G204gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT5), .B(G176gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n314_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT13), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n318_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n318_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(KEYINPUT13), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n303_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n329_), .A2(KEYINPUT72), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(KEYINPUT72), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n285_), .A2(new_n237_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G229gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT73), .ZN(new_n335_));
  INV_X1    g134(.A(new_n285_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n333_), .B(new_n335_), .C1(new_n250_), .C2(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n285_), .A2(new_n237_), .ZN(new_n338_));
  OAI211_X1 g137(.A(G229gat), .B(G233gat), .C1(new_n338_), .C2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G141gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G169gat), .B(G197gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n337_), .A2(new_n339_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n350_));
  OAI22_X1  g149(.A1(new_n350_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(KEYINPUT3), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G141gat), .ZN(new_n357_));
  INV_X1    g156(.A(G148gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n350_), .A3(KEYINPUT3), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n353_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G155gat), .B(G162gat), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(G155gat), .ZN(new_n364_));
  INV_X1    g163(.A(G162gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT1), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(G155gat), .A3(G162gat), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n366_), .B(new_n368_), .C1(G155gat), .C2(G162gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(G141gat), .B(G148gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(G127gat), .A2(G134gat), .ZN(new_n372_));
  INV_X1    g171(.A(G120gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G113gat), .ZN(new_n374_));
  INV_X1    g173(.A(G113gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G120gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G127gat), .A2(G134gat), .ZN(new_n377_));
  AND4_X1   g176(.A1(new_n372_), .A2(new_n374_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n374_), .A2(new_n376_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n363_), .A2(new_n371_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n363_), .B2(new_n371_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n383_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n349_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n363_), .A2(new_n371_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n380_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n361_), .A2(new_n362_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n380_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n349_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n387_), .A2(new_n392_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n392_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(KEYINPUT4), .A3(new_n397_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n348_), .B1(new_n402_), .B2(new_n385_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n403_), .B2(new_n398_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G228gat), .A2(G233gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n407_), .B(KEYINPUT80), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n396_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n412_));
  INV_X1    g211(.A(G218gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n274_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G211gat), .A2(G218gat), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n412_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT21), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G197gat), .B(G204gat), .ZN(new_n418_));
  OR3_X1    g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G197gat), .B(G204gat), .Z(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT21), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n417_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n416_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n409_), .B1(new_n411_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G78gat), .B(G106gat), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n423_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n427_), .B(new_n408_), .C1(new_n396_), .C2(new_n410_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n426_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G22gat), .B(G50gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n393_), .B2(KEYINPUT29), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT79), .B(KEYINPUT28), .ZN(new_n434_));
  INV_X1    g233(.A(new_n432_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n396_), .A2(new_n410_), .A3(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n430_), .A2(new_n431_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n431_), .A2(KEYINPUT82), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441_));
  AOI211_X1 g240(.A(new_n441_), .B(new_n426_), .C1(new_n425_), .C2(new_n428_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n429_), .A2(KEYINPUT83), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n437_), .A2(new_n438_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n425_), .A2(new_n446_), .A3(new_n426_), .A4(new_n428_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n439_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT25), .B(G183gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT26), .B(G190gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT24), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(G169gat), .B2(G176gat), .ZN(new_n456_));
  INV_X1    g255(.A(G169gat), .ZN(new_n457_));
  INV_X1    g256(.A(G176gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n453_), .A2(new_n454_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT23), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(G183gat), .A3(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G183gat), .A2(G190gat), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n463_), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT74), .B1(new_n463_), .B2(KEYINPUT23), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n462_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n460_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(KEYINPUT23), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n462_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G183gat), .A2(G190gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n470_), .A2(new_n472_), .B1(G169gat), .B2(G176gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT22), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G169gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT75), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT22), .B(G169gat), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n458_), .B(new_n476_), .C1(new_n477_), .C2(KEYINPUT75), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n468_), .A2(new_n479_), .A3(KEYINPUT76), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT76), .B1(new_n468_), .B2(new_n479_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n427_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n458_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G169gat), .A2(G176gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n472_), .B2(new_n466_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n460_), .A2(new_n470_), .A3(new_n467_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n427_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT20), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n452_), .B1(new_n482_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G64gat), .B(G92gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G8gat), .B(G36gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n427_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n460_), .A2(new_n470_), .A3(new_n467_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n462_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT74), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n469_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n463_), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n503_), .A2(new_n471_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n498_), .B1(new_n504_), .B2(new_n485_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n505_), .A2(new_n427_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n452_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n497_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n490_), .A2(new_n496_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n470_), .A2(new_n472_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n484_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n476_), .A2(new_n458_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n457_), .A2(KEYINPUT22), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT75), .B1(new_n475_), .B2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n517_));
  AND2_X1   g316(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n518_));
  AND2_X1   g317(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n520_));
  OAI22_X1  g319(.A1(new_n517_), .A2(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n456_), .A2(new_n459_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n467_), .ZN(new_n523_));
  OAI22_X1  g322(.A1(new_n512_), .A2(new_n516_), .B1(new_n523_), .B2(new_n503_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT76), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n468_), .A2(new_n479_), .A3(KEYINPUT76), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n424_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n452_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n507_), .B1(new_n505_), .B2(new_n427_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n532_));
  NAND3_X1  g331(.A1(new_n497_), .A2(new_n506_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n452_), .B2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(KEYINPUT27), .B(new_n510_), .C1(new_n534_), .C2(new_n496_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT27), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n497_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n529_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n495_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n496_), .B1(new_n490_), .B2(new_n509_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n536_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AND4_X1   g340(.A1(new_n406_), .A2(new_n449_), .A3(new_n535_), .A4(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n449_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n539_), .A2(new_n540_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n395_), .A2(KEYINPUT87), .A3(new_n397_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n349_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n392_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n402_), .A2(new_n348_), .A3(new_n385_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(KEYINPUT88), .A3(new_n392_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n392_), .B1(new_n387_), .B2(new_n399_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT33), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n404_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n544_), .A2(new_n554_), .A3(new_n556_), .A4(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n496_), .A2(KEYINPUT32), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n490_), .A2(new_n509_), .A3(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n403_), .A2(new_n401_), .A3(new_n398_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n555_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n531_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n533_), .A2(new_n452_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n560_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT90), .B1(new_n563_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n565_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n560_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT90), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n570_), .A2(new_n405_), .A3(new_n571_), .A4(new_n561_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n559_), .A2(new_n567_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n542_), .B1(new_n543_), .B2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT30), .B(G43gat), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G71gat), .B(G99gat), .Z(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n577_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n526_), .A2(new_n527_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G227gat), .A2(G233gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(G15gat), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n578_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n576_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n578_), .A2(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n582_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n578_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n575_), .A3(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n590_), .A3(KEYINPUT77), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT31), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT31), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n586_), .A2(new_n590_), .A3(KEYINPUT77), .A4(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n394_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n380_), .A3(new_n594_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n592_), .A2(new_n380_), .A3(new_n594_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n380_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n543_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n535_), .A2(new_n541_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT91), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n535_), .A2(new_n541_), .A3(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n406_), .A3(new_n605_), .ZN(new_n606_));
  OAI22_X1  g405(.A1(new_n574_), .A2(new_n598_), .B1(new_n601_), .B2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n330_), .A2(new_n331_), .A3(new_n347_), .A4(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n608_), .A2(G1gat), .A3(new_n406_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT38), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(KEYINPUT38), .ZN(new_n611_));
  INV_X1    g410(.A(new_n347_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n326_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT92), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n267_), .B(KEYINPUT93), .Z(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n302_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n607_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n406_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT94), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n610_), .A2(new_n611_), .A3(new_n619_), .ZN(G1324gat));
  NAND2_X1  g419(.A1(new_n603_), .A2(new_n605_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n608_), .A2(G8gat), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G8gat), .B1(new_n617_), .B2(new_n622_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT96), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT95), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n624_), .B(new_n631_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1325gat));
  NOR2_X1   g434(.A1(new_n599_), .A2(new_n600_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n608_), .A2(G15gat), .A3(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G15gat), .B1(new_n617_), .B2(new_n636_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT41), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1326gat));
  OAI21_X1  g439(.A(G22gat), .B1(new_n617_), .B2(new_n543_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT99), .Z(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT98), .B(KEYINPUT42), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n643_), .ZN(new_n645_));
  OR3_X1    g444(.A1(new_n608_), .A2(G22gat), .A3(new_n543_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n267_), .A2(new_n301_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n613_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(new_n607_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n651_), .A2(G29gat), .A3(new_n406_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n573_), .A2(new_n543_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n542_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n636_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n603_), .A2(new_n406_), .A3(new_n605_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n598_), .A3(new_n543_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n271_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n653_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n607_), .A2(new_n272_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(KEYINPUT101), .A3(new_n661_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n607_), .A2(new_n272_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT102), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n607_), .A2(new_n272_), .A3(new_n669_), .A4(new_n666_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n663_), .A2(new_n665_), .A3(new_n668_), .A4(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n614_), .A2(new_n302_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(KEYINPUT103), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT103), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n671_), .A2(new_n672_), .A3(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n677_), .A3(new_n405_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n652_), .B1(new_n678_), .B2(G29gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT104), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n675_), .A2(new_n677_), .A3(new_n621_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n650_), .A2(new_n683_), .A3(new_n621_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT45), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT105), .B1(new_n682_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1329gat));
  INV_X1    g487(.A(G43gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n650_), .A2(new_n689_), .A3(new_n598_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n675_), .A2(new_n677_), .A3(new_n598_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n689_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT107), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n692_), .B(new_n694_), .ZN(G1330gat));
  OR3_X1    g494(.A1(new_n651_), .A2(G50gat), .A3(new_n543_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n675_), .A2(new_n677_), .A3(new_n449_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n697_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT108), .B1(new_n697_), .B2(G50gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n698_), .B2(new_n699_), .ZN(G1331gat));
  AND3_X1   g499(.A1(new_n607_), .A2(new_n326_), .A3(new_n612_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n616_), .ZN(new_n702_));
  INV_X1    g501(.A(G57gat), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n406_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n303_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(KEYINPUT109), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(KEYINPUT109), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n405_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n704_), .B1(new_n709_), .B2(new_n703_), .ZN(G1332gat));
  OAI21_X1  g509(.A(G64gat), .B1(new_n702_), .B2(new_n622_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n622_), .A2(G64gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n705_), .B2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n702_), .B2(new_n636_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n636_), .A2(G71gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n705_), .B2(new_n717_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n702_), .B2(new_n543_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n543_), .A2(G78gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n705_), .B2(new_n721_), .ZN(G1335gat));
  NAND2_X1  g521(.A1(new_n701_), .A2(new_n648_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT110), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n405_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n327_), .A2(new_n301_), .A3(new_n347_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n671_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n405_), .A2(G85gat), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT111), .Z(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n727_), .B2(new_n729_), .ZN(G1336gat));
  AOI21_X1  g529(.A(G92gat), .B1(new_n724_), .B2(new_n621_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n621_), .A2(new_n226_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n727_), .B2(new_n732_), .ZN(G1337gat));
  AOI21_X1  g532(.A(new_n207_), .B1(new_n727_), .B2(new_n598_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n636_), .A2(new_n222_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n724_), .B2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g536(.A1(new_n671_), .A2(new_n449_), .A3(new_n726_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n671_), .A2(KEYINPUT112), .A3(new_n449_), .A4(new_n726_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n740_), .A2(new_n741_), .A3(G106gat), .A4(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT113), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(G106gat), .A3(new_n742_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT52), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n208_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n741_), .A4(new_n742_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n744_), .A2(new_n746_), .A3(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n724_), .A2(new_n208_), .A3(new_n449_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n750_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1339gat));
  OAI21_X1  g554(.A(KEYINPUT54), .B1(new_n328_), .B2(new_n347_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n303_), .A2(new_n757_), .A3(new_n327_), .A4(new_n612_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n322_), .A2(new_n347_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n307_), .B1(new_n305_), .B2(new_n310_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT55), .ZN(new_n764_));
  INV_X1    g563(.A(new_n311_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n305_), .A2(new_n310_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT55), .A3(new_n306_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n762_), .B(new_n318_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n761_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n311_), .B1(KEYINPUT55), .B2(new_n763_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n768_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n323_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n762_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT56), .B(new_n323_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT115), .A3(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n335_), .B1(new_n338_), .B2(new_n332_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n333_), .B1(new_n250_), .B2(new_n336_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n778_), .B(new_n343_), .C1(new_n779_), .C2(new_n335_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n346_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT116), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n346_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n771_), .A2(new_n777_), .B1(new_n319_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n267_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n775_), .A2(new_n776_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n322_), .A2(new_n785_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n322_), .A2(new_n785_), .A3(KEYINPUT118), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT58), .B1(new_n789_), .B2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n271_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n789_), .A2(new_n794_), .A3(KEYINPUT58), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n788_), .A2(KEYINPUT57), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n771_), .A2(new_n777_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n319_), .A2(new_n785_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n267_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n799_), .B(new_n804_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n760_), .B(new_n798_), .C1(new_n805_), .C2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n302_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT117), .B1(new_n788_), .B2(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n806_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n760_), .B1(new_n811_), .B2(new_n798_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n759_), .B1(new_n809_), .B2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n621_), .A2(new_n406_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n601_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G113gat), .B1(new_n817_), .B2(new_n347_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n803_), .A2(new_n804_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n798_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT120), .B1(new_n820_), .B2(new_n302_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n822_), .B(new_n301_), .C1(new_n798_), .C2(new_n819_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n756_), .A2(new_n758_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n821_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n816_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT121), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n821_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n820_), .A2(KEYINPUT120), .A3(new_n302_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n759_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n826_), .A4(new_n816_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n828_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n826_), .B1(new_n813_), .B2(new_n816_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n375_), .B1(new_n347_), .B2(KEYINPUT122), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(KEYINPUT122), .B2(new_n375_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n818_), .B1(new_n836_), .B2(new_n838_), .ZN(G1340gat));
  OAI21_X1  g638(.A(new_n373_), .B1(new_n327_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n817_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n373_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n834_), .A2(new_n327_), .A3(new_n835_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n373_), .ZN(G1341gat));
  AOI21_X1  g642(.A(G127gat), .B1(new_n817_), .B2(new_n301_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n301_), .A2(G127gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n836_), .B2(new_n845_), .ZN(G1342gat));
  AOI21_X1  g645(.A(G134gat), .B1(new_n817_), .B2(new_n615_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n272_), .A2(G134gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n836_), .B2(new_n848_), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n813_), .A2(new_n636_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n815_), .A2(new_n543_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n850_), .A2(new_n612_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n357_), .ZN(G1344gat));
  NOR3_X1   g653(.A1(new_n850_), .A2(new_n327_), .A3(new_n852_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT123), .B(G148gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1345gat));
  NOR3_X1   g656(.A1(new_n850_), .A2(new_n302_), .A3(new_n852_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT61), .B(G155gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  NAND4_X1  g659(.A1(new_n813_), .A2(new_n636_), .A3(new_n615_), .A4(new_n851_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n365_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n271_), .A2(new_n365_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n813_), .A2(new_n636_), .A3(new_n851_), .A4(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1347gat));
  NOR3_X1   g666(.A1(new_n601_), .A2(new_n622_), .A3(new_n405_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n831_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869_), .B2(new_n612_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(KEYINPUT62), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(KEYINPUT62), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n347_), .A2(new_n477_), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT125), .Z(new_n874_));
  OAI22_X1  g673(.A1(new_n871_), .A2(new_n872_), .B1(new_n869_), .B2(new_n874_), .ZN(G1348gat));
  INV_X1    g674(.A(new_n869_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G176gat), .B1(new_n876_), .B2(new_n326_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n813_), .A2(new_n543_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n622_), .A2(new_n405_), .ZN(new_n879_));
  AND4_X1   g678(.A1(G176gat), .A2(new_n879_), .A3(new_n326_), .A4(new_n598_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n877_), .B1(new_n878_), .B2(new_n880_), .ZN(G1349gat));
  NOR3_X1   g680(.A1(new_n869_), .A2(new_n302_), .A3(new_n453_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n878_), .A2(new_n301_), .A3(new_n598_), .A4(new_n879_), .ZN(new_n883_));
  INV_X1    g682(.A(G183gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1350gat));
  OAI21_X1  g684(.A(G190gat), .B1(new_n869_), .B2(new_n271_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n615_), .A2(new_n454_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n869_), .B2(new_n887_), .ZN(G1351gat));
  NOR3_X1   g687(.A1(new_n622_), .A2(new_n405_), .A3(new_n543_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n813_), .A2(new_n636_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n813_), .A2(new_n892_), .A3(new_n636_), .A4(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G197gat), .B1(new_n894_), .B2(new_n347_), .ZN(new_n895_));
  INV_X1    g694(.A(G197gat), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n896_), .B(new_n612_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1352gat));
  XNOR2_X1  g697(.A(KEYINPUT127), .B(G204gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n894_), .B2(new_n326_), .ZN(new_n901_));
  AOI211_X1 g700(.A(new_n327_), .B(new_n899_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1353gat));
  OR2_X1    g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n894_), .B2(new_n301_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT63), .B(G211gat), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n302_), .B(new_n906_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1354gat));
  NAND2_X1  g707(.A1(new_n894_), .A2(new_n615_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n271_), .A2(new_n413_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n909_), .A2(new_n413_), .B1(new_n894_), .B2(new_n910_), .ZN(G1355gat));
endmodule


