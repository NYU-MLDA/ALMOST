//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G85gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT82), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n211_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n212_), .A2(new_n216_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n207_), .B1(new_n209_), .B2(KEYINPUT1), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n227_), .A2(new_n228_), .B1(new_n229_), .B2(new_n208_), .ZN(new_n230_));
  OAI211_X1 g029(.A(KEYINPUT80), .B(new_n207_), .C1(new_n209_), .C2(KEYINPUT1), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n226_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n224_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT93), .ZN(new_n234_));
  INV_X1    g033(.A(G127gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(G134gat), .ZN(new_n236_));
  INV_X1    g035(.A(G134gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(G127gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT77), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(G127gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(G134gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n242_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n233_), .A2(new_n234_), .A3(new_n245_), .A4(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G155gat), .ZN(new_n251_));
  INV_X1    g050(.A(G162gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT1), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n228_), .B1(new_n253_), .B2(new_n208_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n208_), .A2(new_n229_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n231_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n225_), .ZN(new_n257_));
  INV_X1    g056(.A(G141gat), .ZN(new_n258_));
  INV_X1    g057(.A(G148gat), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n258_), .A2(new_n259_), .B1(KEYINPUT81), .B2(KEYINPUT2), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n219_), .B(new_n218_), .C1(new_n260_), .C2(new_n213_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT82), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n222_), .B(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n210_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n249_), .A2(new_n245_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT93), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n250_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT92), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n257_), .A2(KEYINPUT83), .A3(new_n264_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT83), .B1(new_n257_), .B2(new_n264_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n249_), .A2(KEYINPUT78), .A3(new_n245_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT78), .B1(new_n249_), .B2(new_n245_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n269_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n224_), .B2(new_n232_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n257_), .A2(KEYINPUT83), .A3(new_n264_), .ZN(new_n279_));
  AND4_X1   g078(.A1(new_n269_), .A2(new_n275_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(KEYINPUT4), .B(new_n268_), .C1(new_n276_), .C2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n272_), .A2(new_n282_), .A3(new_n275_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G225gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n268_), .B(new_n284_), .C1(new_n276_), .C2(new_n280_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n206_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n206_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n250_), .A2(new_n267_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n249_), .A2(new_n245_), .A3(KEYINPUT78), .ZN(new_n293_));
  INV_X1    g092(.A(new_n274_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n278_), .A2(new_n293_), .A3(new_n294_), .A4(new_n279_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT92), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n275_), .A2(new_n269_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n292_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n286_), .B1(new_n298_), .B2(KEYINPUT4), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT96), .B1(new_n291_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n206_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n298_), .B2(new_n284_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT96), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n288_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n290_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G183gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT25), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT25), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G183gat), .ZN(new_n309_));
  INV_X1    g108(.A(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT26), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G190gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n307_), .A2(new_n309_), .A3(new_n311_), .A4(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT23), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(G183gat), .A3(G190gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(KEYINPUT72), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(G169gat), .B2(G176gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326_));
  AND4_X1   g125(.A1(KEYINPUT24), .A2(new_n323_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT24), .B1(new_n323_), .B2(new_n325_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n320_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n326_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n319_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n315_), .B2(KEYINPUT23), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n306_), .A2(new_n310_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n330_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n321_), .B2(KEYINPUT22), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT73), .A3(G169gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n321_), .A2(KEYINPUT22), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n339_), .A2(new_n341_), .A3(new_n322_), .A4(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT74), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n329_), .B1(new_n337_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(G197gat), .B(G204gat), .Z(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(KEYINPUT85), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G197gat), .B(G204gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT21), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT21), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT90), .B1(new_n345_), .B2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n354_), .B2(new_n348_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n343_), .B(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n333_), .B1(new_n319_), .B2(new_n331_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n336_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n326_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n328_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(new_n319_), .A3(new_n314_), .ZN(new_n366_));
  OAI22_X1  g165(.A1(new_n361_), .A2(new_n364_), .B1(new_n327_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT90), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n359_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n357_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT19), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT20), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n340_), .A2(G169gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n342_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n326_), .B1(new_n376_), .B2(G176gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n319_), .A2(new_n336_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT89), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT89), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n319_), .A2(new_n380_), .A3(new_n336_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n377_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n326_), .A2(new_n383_), .A3(KEYINPUT24), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n326_), .B2(KEYINPUT24), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n314_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT88), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT88), .B(new_n314_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n362_), .A2(new_n328_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n382_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n374_), .B1(new_n393_), .B2(new_n356_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n370_), .A2(new_n373_), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n393_), .A2(new_n356_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT20), .B1(new_n359_), .B2(new_n367_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n372_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT18), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n399_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT95), .ZN(new_n408_));
  INV_X1    g207(.A(new_n397_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n409_), .B(new_n373_), .C1(new_n356_), .C2(new_n393_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n390_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n326_), .A2(KEYINPUT24), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT87), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n413_), .A2(new_n323_), .A3(new_n325_), .A4(new_n384_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT88), .B1(new_n414_), .B2(new_n314_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n392_), .B1(new_n411_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n382_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n356_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT20), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n357_), .B2(new_n369_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n410_), .B1(new_n420_), .B2(new_n373_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n408_), .B1(new_n421_), .B2(new_n405_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n373_), .B1(new_n370_), .B2(new_n394_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n396_), .A2(new_n397_), .A3(new_n372_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n408_), .B(new_n405_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n407_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n202_), .B1(new_n305_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n289_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n301_), .B1(new_n299_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n288_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n303_), .B1(new_n288_), .B2(new_n302_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n405_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT95), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n406_), .B1(new_n435_), .B2(new_n425_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(KEYINPUT97), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT94), .B1(new_n291_), .B2(new_n299_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT94), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n288_), .A2(new_n302_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n399_), .A2(new_n403_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n395_), .A2(new_n398_), .A3(new_n404_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT91), .A3(new_n444_), .ZN(new_n445_));
  OR3_X1    g244(.A1(new_n399_), .A2(KEYINPUT91), .A3(new_n403_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n288_), .A2(new_n302_), .A3(KEYINPUT33), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n281_), .A2(new_n284_), .A3(new_n283_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n206_), .B1(new_n298_), .B2(new_n285_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n442_), .A2(new_n447_), .A3(new_n448_), .A4(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n428_), .A2(new_n437_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n278_), .A2(new_n279_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT28), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT29), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n455_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT84), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n457_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G22gat), .B(G50gat), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n460_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n356_), .B1(G228gat), .B2(G233gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n456_), .B2(new_n454_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n472_));
  OAI21_X1  g271(.A(new_n359_), .B1(new_n233_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(G228gat), .A3(G233gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G78gat), .B(G106gat), .Z(new_n476_));
  AND2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n475_), .A2(new_n476_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n469_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n453_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n305_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n445_), .A2(new_n446_), .A3(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n423_), .A2(new_n424_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(new_n404_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n444_), .A2(KEYINPUT27), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT98), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n421_), .A2(new_n403_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT98), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(KEYINPUT27), .A4(new_n444_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n487_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n485_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n484_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT100), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n275_), .B(KEYINPUT79), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(KEYINPUT31), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(KEYINPUT31), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT76), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G227gat), .A2(G233gat), .ZN(new_n504_));
  INV_X1    g303(.A(G15gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT30), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n503_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G43gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n367_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n508_), .B(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n498_), .A2(new_n499_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n496_), .B1(new_n453_), .B2(new_n483_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n512_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT100), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n495_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n515_), .A2(new_n483_), .A3(new_n305_), .A4(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT12), .ZN(new_n520_));
  XOR2_X1   g319(.A(G85gat), .B(G92gat), .Z(new_n521_));
  INV_X1    g320(.A(KEYINPUT8), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT6), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(G99gat), .A3(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT64), .ZN(new_n529_));
  NOR2_X1   g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT7), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n523_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n528_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n522_), .B1(new_n533_), .B2(new_n521_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT10), .B(G99gat), .Z(new_n536_));
  INV_X1    g335(.A(G106gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT9), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(G85gat), .A3(G92gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n521_), .A2(KEYINPUT9), .ZN(new_n541_));
  AND4_X1   g340(.A1(new_n529_), .A2(new_n538_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT11), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT65), .ZN(new_n546_));
  XOR2_X1   g345(.A(G71gat), .B(G78gat), .Z(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(KEYINPUT11), .B2(new_n544_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n546_), .B(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n520_), .B1(new_n543_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n549_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n543_), .A2(KEYINPUT66), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT66), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n535_), .B2(new_n542_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n549_), .A2(new_n520_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n552_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n553_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n551_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n543_), .A2(new_n549_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT67), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n559_), .A2(new_n563_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT13), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n570_), .A2(KEYINPUT13), .A3(new_n572_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578_));
  INV_X1    g377(.A(G1gat), .ZN(new_n579_));
  INV_X1    g378(.A(G8gat), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT14), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G1gat), .B(G8gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G29gat), .B(G36gat), .Z(new_n585_));
  XOR2_X1   g384(.A(G43gat), .B(G50gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n584_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT69), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n587_), .B(KEYINPUT15), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n584_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n584_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n587_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(new_n590_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n589_), .A2(new_n591_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT71), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT70), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n597_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n577_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n519_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n554_), .A2(new_n592_), .A3(new_n556_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT35), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT34), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n543_), .A2(new_n587_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n612_), .A2(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n614_), .A2(new_n615_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n622_), .B(KEYINPUT36), .Z(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT37), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n627_), .A2(KEYINPUT37), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(G127gat), .B(G155gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT16), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT68), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(new_n584_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(new_n549_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(new_n636_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n549_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n631_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n607_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n579_), .A3(new_n433_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n519_), .A2(new_n645_), .A3(new_n627_), .A4(new_n606_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n305_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n650_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n653_), .A3(new_n654_), .ZN(G1324gat));
  OAI21_X1  g454(.A(G8gat), .B1(new_n652_), .B2(new_n517_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT39), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n648_), .A2(new_n580_), .A3(new_n495_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g459(.A(G15gat), .B1(new_n652_), .B2(new_n512_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT41), .Z(new_n662_));
  NAND3_X1  g461(.A1(new_n648_), .A2(new_n505_), .A3(new_n515_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  OAI21_X1  g463(.A(G22gat), .B1(new_n652_), .B2(new_n483_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n483_), .A2(G22gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n647_), .B2(new_n667_), .ZN(G1327gat));
  NOR2_X1   g467(.A1(new_n645_), .A2(new_n627_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n607_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n433_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n631_), .A2(KEYINPUT43), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n519_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n519_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n513_), .A2(new_n516_), .A3(KEYINPUT101), .A4(new_n518_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n631_), .B(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(new_n677_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n674_), .B1(new_n681_), .B2(KEYINPUT43), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n606_), .A2(new_n644_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n672_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n683_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n679_), .B1(new_n519_), .B2(new_n675_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(new_n677_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n685_), .C1(new_n688_), .C2(new_n674_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n684_), .A2(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n433_), .A2(G29gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n671_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n495_), .A3(new_n689_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n517_), .A2(G36gat), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n670_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT104), .Z(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n670_), .A2(new_n696_), .A3(new_n699_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n695_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n693_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n703_), .B1(new_n694_), .B2(G36gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n708_), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710_));
  AND4_X1   g509(.A1(new_n710_), .A2(new_n695_), .A3(KEYINPUT46), .A4(new_n704_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n708_), .B2(KEYINPUT46), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n707_), .A2(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1329gat));
  INV_X1    g512(.A(G43gat), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n512_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n684_), .A2(new_n689_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n684_), .A2(new_n689_), .A3(KEYINPUT107), .A4(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n670_), .A2(new_n515_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n714_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g522(.A(G50gat), .ZN(new_n724_));
  INV_X1    g523(.A(new_n483_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n670_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n690_), .A2(KEYINPUT108), .A3(new_n725_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G50gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT108), .B1(new_n690_), .B2(new_n725_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(G1331gat));
  INV_X1    g529(.A(new_n577_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n604_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n519_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n646_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n433_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT109), .Z(new_n736_));
  NAND4_X1  g535(.A1(new_n519_), .A2(new_n645_), .A3(new_n627_), .A4(new_n732_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT110), .Z(new_n738_));
  AND2_X1   g537(.A1(new_n433_), .A2(G57gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n495_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G64gat), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT48), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n517_), .A2(G64gat), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT111), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n734_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(G1333gat));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n734_), .A2(new_n748_), .A3(new_n515_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n738_), .A2(new_n515_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G71gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT49), .B(new_n748_), .C1(new_n738_), .C2(new_n515_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(G1334gat));
  INV_X1    g555(.A(G78gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n738_), .B2(new_n725_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT50), .Z(new_n759_));
  NAND3_X1  g558(.A1(new_n734_), .A2(new_n757_), .A3(new_n725_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1335gat));
  INV_X1    g560(.A(new_n682_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n732_), .A2(new_n644_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n305_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n733_), .A2(new_n669_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n305_), .A2(G85gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n765_), .B2(new_n517_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n517_), .A2(G92gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n767_), .B2(new_n771_), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n765_), .B2(new_n512_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n767_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n536_), .A3(new_n515_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n537_), .A3(new_n725_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n762_), .A2(new_n725_), .A3(new_n764_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n778_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NOR4_X1   g586(.A1(new_n512_), .A2(new_n725_), .A3(new_n305_), .A4(new_n495_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT120), .Z(new_n789_));
  INV_X1    g588(.A(new_n627_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n570_), .A2(new_n791_), .A3(new_n604_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n570_), .B2(new_n604_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n559_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n559_), .B2(new_n795_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n553_), .B1(new_n552_), .B2(new_n558_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT116), .B1(new_n800_), .B2(new_n568_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n559_), .A2(new_n795_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT55), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n559_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n799_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n567_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .A4(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n798_), .A2(new_n799_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n568_), .B1(new_n812_), .B2(new_n806_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n808_), .A2(new_n567_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT56), .B1(new_n816_), .B2(KEYINPUT116), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n802_), .B1(new_n817_), .B2(new_n810_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n794_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n589_), .A2(new_n590_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT118), .B1(new_n820_), .B2(new_n602_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n590_), .B1(new_n594_), .B2(new_n587_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n593_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(KEYINPUT118), .A3(new_n602_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n823_), .A2(new_n824_), .B1(new_n601_), .B2(new_n597_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n573_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n790_), .B1(new_n819_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT119), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n570_), .A2(new_n825_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n816_), .A2(new_n803_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n814_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT58), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(KEYINPUT58), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n631_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n827_), .A2(new_n829_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n803_), .B1(new_n813_), .B2(new_n809_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n810_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT117), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n814_), .A3(new_n811_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n840_), .A2(new_n794_), .B1(new_n573_), .B2(new_n825_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT119), .B(new_n828_), .C1(new_n841_), .C2(new_n790_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n645_), .B1(new_n836_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n644_), .A2(new_n604_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT113), .B1(new_n731_), .B2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n575_), .A2(KEYINPUT113), .A3(new_n576_), .A4(new_n844_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n631_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT54), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n789_), .B1(new_n843_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n604_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT121), .B1(new_n843_), .B2(new_n849_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n850_), .A3(new_n855_), .ZN(new_n856_));
  OAI221_X1 g655(.A(new_n789_), .B1(KEYINPUT121), .B2(KEYINPUT59), .C1(new_n843_), .C2(new_n849_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n605_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n853_), .B1(new_n858_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860_));
  AOI21_X1  g659(.A(G120gat), .B1(new_n577_), .B2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n860_), .B2(G120gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n851_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n731_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n864_));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT122), .B(new_n863_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1341gat));
  AOI21_X1  g669(.A(G127gat), .B1(new_n851_), .B2(new_n645_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n856_), .A2(new_n857_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n645_), .A2(G127gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT123), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n871_), .B1(new_n872_), .B2(new_n874_), .ZN(G1342gat));
  NOR2_X1   g674(.A1(new_n631_), .A2(new_n237_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G134gat), .B1(new_n851_), .B2(new_n790_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT124), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n878_), .A2(new_n880_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n843_), .A2(new_n849_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n512_), .A2(new_n725_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n495_), .A2(new_n305_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n888_), .A2(KEYINPUT125), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT125), .B1(new_n888_), .B2(new_n889_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n604_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G141gat), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n258_), .B(new_n604_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1344gat));
  OAI21_X1  g694(.A(new_n577_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G148gat), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n259_), .B(new_n577_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1345gat));
  OAI21_X1  g698(.A(new_n645_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n901_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n645_), .B(new_n903_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1346gat));
  OR2_X1    g704(.A1(new_n890_), .A2(new_n891_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n679_), .A2(new_n252_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n790_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n906_), .A2(new_n907_), .B1(new_n908_), .B2(new_n252_), .ZN(G1347gat));
  OR2_X1    g708(.A1(new_n843_), .A2(new_n849_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n512_), .A2(new_n517_), .A3(new_n725_), .A4(new_n433_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT126), .B1(new_n912_), .B2(new_n605_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n910_), .A2(new_n914_), .A3(new_n604_), .A4(new_n911_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(G169gat), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n913_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n915_), .ZN(new_n919_));
  OR3_X1    g718(.A1(new_n912_), .A2(new_n376_), .A3(new_n605_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(G1348gat));
  NOR2_X1   g720(.A1(new_n912_), .A2(new_n731_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n322_), .ZN(G1349gat));
  NOR2_X1   g722(.A1(new_n912_), .A2(new_n644_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(G183gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n307_), .A2(new_n309_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n924_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n912_), .B2(new_n631_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n790_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n912_), .B2(new_n929_), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n517_), .A2(new_n433_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n888_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n604_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n577_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g736(.A1(new_n932_), .A2(new_n644_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AND2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n938_), .B2(new_n939_), .ZN(G1354gat));
  AOI21_X1  g741(.A(G218gat), .B1(new_n933_), .B2(new_n790_), .ZN(new_n943_));
  INV_X1    g742(.A(G218gat), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n631_), .A2(new_n944_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT127), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n943_), .B1(new_n933_), .B2(new_n946_), .ZN(G1355gat));
endmodule


