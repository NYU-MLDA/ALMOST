//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(G15gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT76), .B(G176gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT22), .B(G169gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT77), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n212_), .A2(KEYINPUT78), .A3(G183gat), .A4(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT23), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI221_X1 g017(.A(new_n213_), .B1(G183gat), .B2(G190gat), .C1(new_n218_), .C2(KEYINPUT78), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n208_), .A2(new_n220_), .A3(new_n209_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n211_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G169gat), .ZN(new_n226_));
  INV_X1    g025(.A(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(KEYINPUT24), .A3(new_n209_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(KEYINPUT24), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n225_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n218_), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n222_), .A2(KEYINPUT79), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT79), .B1(new_n222_), .B2(new_n232_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n205_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n222_), .A2(new_n232_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n222_), .A2(KEYINPUT79), .A3(new_n232_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n205_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G71gat), .B(G99gat), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n235_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n202_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n235_), .A2(new_n241_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n245_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n235_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(KEYINPUT82), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT81), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n248_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n202_), .B(new_n260_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT83), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT3), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  AND2_X1   g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n274_), .A2(new_n276_), .B1(KEYINPUT2), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n272_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT86), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT86), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n278_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n269_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n267_), .B1(KEYINPUT1), .B2(new_n268_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT84), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT84), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n284_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n288_), .A2(new_n277_), .A3(new_n273_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n283_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n291_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G22gat), .B(G50gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n283_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n289_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n292_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT28), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n296_), .B1(new_n302_), .B2(new_n293_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n265_), .B1(new_n298_), .B2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(G228gat), .A2(G233gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(KEYINPUT87), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT29), .B1(new_n283_), .B2(new_n289_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G197gat), .B(G204gat), .Z(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n306_), .B1(new_n307_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G78gat), .B(G106gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n305_), .A2(KEYINPUT87), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  AOI211_X1 g119(.A(new_n306_), .B(new_n318_), .C1(new_n307_), .C2(new_n314_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n297_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n302_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(KEYINPUT88), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n304_), .A2(new_n323_), .A3(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n322_), .A2(KEYINPUT88), .A3(new_n325_), .A4(new_n324_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n259_), .A2(KEYINPUT83), .A3(new_n261_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n264_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n329_), .B2(new_n262_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT27), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT20), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n233_), .A2(new_n234_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n314_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341_));
  MUX2_X1   g140(.A(new_n217_), .B(new_n218_), .S(new_n341_), .Z(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n231_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n210_), .A2(KEYINPUT89), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n210_), .B2(KEYINPUT89), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n343_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n314_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT90), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT90), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n350_), .A3(new_n314_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n336_), .B1(new_n340_), .B2(new_n352_), .ZN(new_n353_));
  OR3_X1    g152(.A1(new_n347_), .A2(KEYINPUT91), .A3(new_n314_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT91), .B1(new_n347_), .B2(new_n314_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n238_), .A2(new_n239_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n314_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n335_), .A2(new_n337_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT18), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n353_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n352_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n357_), .B2(new_n314_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n335_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n364_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n333_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n367_), .A2(new_n368_), .A3(new_n335_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n357_), .B2(new_n314_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT96), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n314_), .B1(new_n347_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n376_), .B2(new_n347_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n336_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n365_), .B1(new_n373_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n369_), .A2(new_n364_), .A3(new_n370_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(KEYINPUT27), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n372_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n257_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n290_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n257_), .B1(new_n283_), .B2(new_n289_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(KEYINPUT4), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n387_), .A2(KEYINPUT4), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n384_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G1gat), .B(G29gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT92), .B(G85gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  INV_X1    g194(.A(new_n384_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n397_));
  OR3_X1    g196(.A1(new_n390_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(new_n390_), .B2(new_n397_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n383_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n369_), .A2(new_n370_), .A3(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT32), .B(new_n364_), .C1(new_n373_), .C2(new_n379_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n371_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT33), .B(new_n395_), .C1(new_n390_), .C2(new_n397_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n388_), .A2(new_n384_), .A3(new_n389_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n395_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n386_), .A2(new_n396_), .A3(new_n387_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n406_), .A2(new_n381_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n399_), .A2(KEYINPUT93), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT93), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n415_), .B(new_n395_), .C1(new_n390_), .C2(new_n397_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n413_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n405_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n259_), .A2(KEYINPUT83), .A3(new_n261_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT83), .B1(new_n259_), .B2(new_n261_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n419_), .A2(new_n329_), .A3(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n332_), .A2(new_n401_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G190gat), .B(G218gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G134gat), .B(G162gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT36), .Z(new_n426_));
  XNOR2_X1  g225(.A(G29gat), .B(G36gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT67), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G43gat), .B(G50gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT67), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n427_), .B(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT10), .B(G99gat), .Z(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G85gat), .A2(G92gat), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n439_), .A2(KEYINPUT9), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G99gat), .A2(G106gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(KEYINPUT9), .A3(new_n439_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n438_), .A2(new_n440_), .A3(new_n445_), .A4(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  INV_X1    g248(.A(G99gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n437_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n451_), .A2(new_n443_), .A3(new_n444_), .A4(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT8), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n446_), .A2(new_n439_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n448_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G232gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT34), .ZN(new_n460_));
  OAI22_X1  g259(.A1(new_n435_), .A2(new_n458_), .B1(KEYINPUT35), .B2(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n430_), .A2(new_n434_), .A3(KEYINPUT15), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT15), .B1(new_n430_), .B2(new_n434_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n464_), .B2(new_n458_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n460_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT35), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n465_), .A2(new_n469_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n426_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n472_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n425_), .A2(KEYINPUT36), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n422_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G127gat), .B(G155gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT16), .ZN(new_n481_));
  XOR2_X1   g280(.A(G183gat), .B(G211gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT17), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G1gat), .B(G8gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT70), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  INV_X1    g288(.A(G1gat), .ZN(new_n490_));
  INV_X1    g289(.A(G8gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n486_), .B(KEYINPUT70), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G231gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G57gat), .B(G64gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G71gat), .B(G78gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT11), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(KEYINPUT11), .ZN(new_n504_));
  INV_X1    g303(.A(new_n502_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n501_), .A2(KEYINPUT11), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n503_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n500_), .B(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(KEYINPUT17), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n485_), .B1(new_n510_), .B2(new_n483_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n509_), .A2(KEYINPUT71), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n453_), .A2(new_n455_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT8), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n508_), .B1(new_n517_), .B2(new_n448_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT65), .B1(new_n518_), .B2(KEYINPUT66), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT12), .B1(new_n518_), .B2(KEYINPUT65), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G230gat), .A2(G233gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n522_), .B(KEYINPUT64), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n458_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n508_), .ZN(new_n526_));
  OAI211_X1 g325(.A(KEYINPUT65), .B(KEYINPUT12), .C1(new_n518_), .C2(KEYINPUT66), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n521_), .A2(new_n524_), .A3(new_n526_), .A4(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n526_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n523_), .B1(new_n529_), .B2(new_n518_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G120gat), .B(G148gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT5), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n528_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n495_), .B(new_n497_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n496_), .A2(new_n493_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n488_), .A2(new_n494_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n430_), .B(new_n434_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n435_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n547_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n548_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT72), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n554_));
  AOI211_X1 g353(.A(new_n554_), .B(new_n548_), .C1(new_n550_), .C2(new_n547_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n549_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n549_), .B(new_n563_), .C1(new_n553_), .C2(new_n555_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n543_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n479_), .A2(new_n513_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n400_), .ZN(new_n569_));
  OAI21_X1  g368(.A(G1gat), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT98), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n565_), .B(KEYINPUT75), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n422_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT69), .B1(new_n477_), .B2(KEYINPUT37), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n473_), .A2(new_n476_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n426_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n474_), .B2(new_n470_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(KEYINPUT68), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n476_), .B1(new_n580_), .B2(KEYINPUT68), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT37), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n513_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n543_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n573_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n573_), .A2(KEYINPUT97), .A3(new_n586_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n589_), .A2(new_n490_), .A3(new_n400_), .A4(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n571_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT99), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n571_), .A2(new_n593_), .A3(new_n597_), .A4(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(G1324gat));
  INV_X1    g398(.A(new_n383_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G8gat), .B1(new_n568_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT39), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n589_), .A2(new_n491_), .A3(new_n383_), .A4(new_n590_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n604_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1325gat));
  NOR2_X1   g407(.A1(new_n419_), .A2(new_n420_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n587_), .A2(G15gat), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT101), .ZN(new_n611_));
  OAI21_X1  g410(.A(G15gat), .B1(new_n568_), .B2(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n613_), .A3(new_n614_), .ZN(G1326gat));
  XNOR2_X1  g414(.A(new_n329_), .B(KEYINPUT102), .ZN(new_n616_));
  OAI21_X1  g415(.A(G22gat), .B1(new_n568_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT42), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n616_), .A2(G22gat), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n618_), .B1(new_n587_), .B2(new_n619_), .ZN(G1327gat));
  INV_X1    g419(.A(new_n513_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT43), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n327_), .A2(new_n328_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n419_), .A2(new_n420_), .A3(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n329_), .A2(new_n262_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n401_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n421_), .A2(new_n418_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n584_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n622_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT43), .B(new_n584_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n621_), .B(new_n567_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT103), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n567_), .A2(new_n621_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT43), .B1(new_n422_), .B2(new_n584_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n622_), .A3(new_n629_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n633_), .A2(new_n634_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n400_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT104), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n633_), .A2(new_n640_), .A3(new_n634_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n400_), .A4(new_n642_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n644_), .A2(G29gat), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n621_), .A2(new_n478_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT105), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n543_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n573_), .ZN(new_n652_));
  OR3_X1    g451(.A1(new_n652_), .A2(G29gat), .A3(new_n569_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n648_), .A2(new_n653_), .ZN(G1328gat));
  NAND2_X1  g453(.A1(new_n642_), .A2(new_n383_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G36gat), .B1(new_n641_), .B2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n383_), .A2(new_n658_), .ZN(new_n659_));
  OR3_X1    g458(.A1(new_n652_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n652_), .B2(new_n659_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n656_), .A2(KEYINPUT46), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(new_n655_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n658_), .B1(new_n666_), .B2(new_n645_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n667_), .B2(new_n662_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(G1329gat));
  XNOR2_X1  g468(.A(KEYINPUT107), .B(G43gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n652_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n609_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n262_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n642_), .A2(G43gat), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n675_), .B2(new_n645_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT47), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1330gat));
  INV_X1    g477(.A(new_n616_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G50gat), .B1(new_n671_), .B2(new_n679_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n642_), .A2(G50gat), .A3(new_n329_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n645_), .ZN(G1331gat));
  INV_X1    g481(.A(new_n543_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n572_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n621_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n479_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G57gat), .B1(new_n686_), .B2(new_n569_), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n422_), .A2(new_n565_), .A3(new_n683_), .A4(new_n585_), .ZN(new_n688_));
  INV_X1    g487(.A(G57gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n400_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(G1332gat));
  OAI21_X1  g490(.A(G64gat), .B1(new_n686_), .B2(new_n600_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n692_), .B(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n696_), .A3(new_n383_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g498(.A(G71gat), .B1(new_n686_), .B2(new_n609_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT49), .ZN(new_n701_));
  INV_X1    g500(.A(G71gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n688_), .A2(new_n702_), .A3(new_n672_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1334gat));
  OAI21_X1  g503(.A(G78gat), .B1(new_n686_), .B2(new_n616_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT50), .ZN(new_n706_));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n688_), .A2(new_n707_), .A3(new_n679_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1335gat));
  INV_X1    g508(.A(G85gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n650_), .A2(new_n683_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n628_), .A3(new_n566_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n712_), .B2(new_n569_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT110), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n636_), .A2(new_n637_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n683_), .A2(new_n565_), .A3(new_n513_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT111), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n400_), .A2(G85gat), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT112), .Z(new_n721_));
  AOI21_X1  g520(.A(new_n714_), .B1(new_n719_), .B2(new_n721_), .ZN(G1336gat));
  OAI21_X1  g521(.A(G92gat), .B1(new_n718_), .B2(new_n600_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n600_), .A2(G92gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n712_), .B2(new_n724_), .ZN(G1337gat));
  NAND2_X1  g524(.A1(new_n674_), .A2(new_n436_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n712_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT113), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n717_), .A2(new_n672_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n728_), .B(new_n729_), .C1(new_n450_), .C2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n727_), .B(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(new_n450_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT51), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n735_), .ZN(G1338gat));
  OR3_X1    g535(.A1(new_n712_), .A2(G106gat), .A3(new_n623_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n329_), .B(new_n716_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n715_), .A2(KEYINPUT114), .A3(new_n329_), .A4(new_n716_), .ZN(new_n742_));
  AND4_X1   g541(.A1(new_n738_), .A2(new_n741_), .A3(G106gat), .A4(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n437_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n738_), .B1(new_n744_), .B2(new_n742_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n737_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n737_), .C1(new_n743_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  NAND4_X1  g549(.A1(new_n683_), .A2(new_n584_), .A3(new_n572_), .A4(new_n513_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n544_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n563_), .B1(new_n551_), .B2(new_n548_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n564_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n536_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT65), .ZN(new_n759_));
  INV_X1    g558(.A(new_n508_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n458_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT66), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT12), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n761_), .B2(new_n759_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n527_), .B(new_n526_), .C1(new_n763_), .C2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n523_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n528_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n529_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n772_), .A2(KEYINPUT55), .A3(new_n524_), .A4(new_n527_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n766_), .A2(KEYINPUT115), .A3(new_n523_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n769_), .A2(new_n771_), .A3(new_n773_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n534_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n534_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n758_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT58), .B1(new_n780_), .B2(KEYINPUT118), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n534_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n534_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n782_), .B(new_n783_), .C1(new_n786_), .C2(new_n758_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n781_), .A2(new_n629_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n757_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT117), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n757_), .B(new_n792_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n778_), .A2(new_n795_), .A3(new_n779_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n775_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n534_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n537_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n794_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n789_), .B1(new_n800_), .B2(new_n478_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n794_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n784_), .A2(new_n785_), .A3(KEYINPUT116), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n798_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n478_), .A2(new_n789_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n788_), .A2(new_n801_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n513_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n788_), .A2(new_n801_), .A3(KEYINPUT119), .A4(new_n807_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n753_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n383_), .A2(new_n569_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n625_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT59), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n808_), .A2(new_n621_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n751_), .B(KEYINPUT54), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n814_), .ZN(new_n819_));
  XOR2_X1   g618(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n820_));
  AND2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n815_), .A2(new_n684_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G113gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n808_), .A2(new_n809_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n621_), .A3(new_n811_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n817_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n819_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n566_), .A2(G113gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n828_), .B2(new_n829_), .ZN(G1340gat));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n831_));
  AOI21_X1  g630(.A(G120gat), .B1(new_n543_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n831_), .B2(G120gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n827_), .A2(new_n819_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n822_), .A2(new_n543_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n828_), .B2(KEYINPUT59), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT121), .B(new_n834_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n683_), .B1(new_n818_), .B2(new_n821_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n837_), .B1(new_n815_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n834_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n839_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n838_), .A2(new_n843_), .ZN(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n828_), .B2(new_n621_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n513_), .B2(KEYINPUT122), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(KEYINPUT122), .B2(new_n845_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n815_), .A2(new_n822_), .A3(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n846_), .A2(new_n849_), .ZN(G1342gat));
  NAND3_X1  g649(.A1(new_n815_), .A2(new_n629_), .A3(new_n822_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G134gat), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n477_), .A2(G134gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n828_), .B2(new_n853_), .ZN(G1343gat));
  NOR2_X1   g653(.A1(new_n812_), .A2(new_n331_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n565_), .A3(new_n813_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT123), .B(G141gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1344gat));
  NAND3_X1  g657(.A1(new_n855_), .A2(new_n543_), .A3(new_n813_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT124), .B(G148gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1345gat));
  NAND3_X1  g660(.A1(new_n855_), .A2(new_n513_), .A3(new_n813_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  AND4_X1   g663(.A1(G162gat), .A2(new_n855_), .A3(new_n629_), .A4(new_n813_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n855_), .A2(new_n478_), .A3(new_n813_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT125), .ZN(new_n867_));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n813_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n812_), .A2(new_n331_), .A3(new_n477_), .A4(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT125), .B1(new_n871_), .B2(G162gat), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n865_), .B1(new_n869_), .B2(new_n872_), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n600_), .A2(new_n400_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n609_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n679_), .B(new_n877_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n226_), .B1(new_n878_), .B2(new_n565_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n879_), .A2(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(KEYINPUT62), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n207_), .A3(new_n565_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  NAND2_X1  g682(.A1(new_n878_), .A2(new_n543_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n812_), .A2(new_n329_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n877_), .A2(new_n227_), .A3(new_n683_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n884_), .A2(new_n206_), .B1(new_n885_), .B2(new_n886_), .ZN(G1349gat));
  NAND3_X1  g686(.A1(new_n885_), .A2(new_n513_), .A3(new_n876_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n621_), .A2(new_n223_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n888_), .A2(new_n214_), .B1(new_n878_), .B2(new_n889_), .ZN(G1350gat));
  AND3_X1   g689(.A1(new_n878_), .A2(new_n224_), .A3(new_n478_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n215_), .B1(new_n878_), .B2(new_n629_), .ZN(new_n892_));
  OR3_X1    g691(.A1(new_n891_), .A2(new_n892_), .A3(KEYINPUT126), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT126), .B1(new_n891_), .B2(new_n892_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1351gat));
  AOI211_X1 g694(.A(new_n331_), .B(new_n875_), .C1(new_n826_), .C2(new_n817_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n565_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n543_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g699(.A(KEYINPUT63), .B(G211gat), .Z(new_n901_));
  AND3_X1   g700(.A1(new_n896_), .A2(new_n513_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n896_), .A2(new_n513_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(G1354gat));
  INV_X1    g704(.A(G218gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n896_), .B2(new_n629_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n477_), .A2(G218gat), .ZN(new_n908_));
  AND4_X1   g707(.A1(new_n624_), .A2(new_n827_), .A3(new_n874_), .A4(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT127), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n896_), .A2(new_n908_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n812_), .A2(new_n331_), .A3(new_n584_), .A4(new_n875_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n911_), .B(new_n912_), .C1(new_n913_), .C2(new_n906_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(G1355gat));
endmodule


