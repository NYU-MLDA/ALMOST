//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT91), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT91), .ZN(new_n204_));
  INV_X1    g003(.A(G211gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(G218gat), .ZN(new_n206_));
  INV_X1    g005(.A(G218gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(G211gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n203_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G197gat), .ZN(new_n211_));
  INV_X1    g010(.A(G204gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT89), .B(G204gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(new_n211_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT92), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(KEYINPUT92), .B(new_n213_), .C1(new_n214_), .C2(new_n211_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n210_), .A2(new_n217_), .A3(KEYINPUT21), .A4(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n214_), .A2(G197gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT88), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(new_n211_), .B2(G204gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n212_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT21), .B1(new_n220_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n215_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n203_), .A2(new_n209_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G183gat), .ZN(new_n233_));
  INV_X1    g032(.A(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT26), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G190gat), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n231_), .A2(new_n233_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(KEYINPUT24), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n238_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(G183gat), .A3(G190gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT80), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT80), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n249_), .A2(new_n246_), .A3(G183gat), .A4(G190gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n248_), .A2(new_n250_), .B1(KEYINPUT23), .B2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(KEYINPUT23), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n247_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(KEYINPUT81), .A2(G169gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT22), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT22), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(KEYINPUT81), .A3(G169gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .A4(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n265_), .A3(new_n241_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n219_), .A2(new_n229_), .A3(new_n253_), .A4(new_n266_), .ZN(new_n267_));
  AND4_X1   g066(.A1(KEYINPUT21), .A2(new_n218_), .A3(new_n203_), .A4(new_n209_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n215_), .A2(new_n226_), .B1(new_n203_), .B2(new_n209_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n268_), .A2(new_n217_), .B1(new_n225_), .B2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n263_), .A2(new_n264_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT22), .B(G169gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n241_), .B(new_n273_), .C1(new_n252_), .C2(new_n256_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n238_), .A2(new_n242_), .A3(new_n244_), .A4(new_n255_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n267_), .B(KEYINPUT20), .C1(new_n270_), .C2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT19), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT94), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G8gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT18), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G64gat), .ZN(new_n286_));
  INV_X1    g085(.A(G92gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n278_), .A2(KEYINPUT94), .A3(new_n280_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n219_), .A2(new_n229_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT20), .B1(new_n290_), .B2(new_n276_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n219_), .A2(new_n229_), .B1(new_n253_), .B2(new_n266_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n280_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n283_), .A2(new_n288_), .A3(new_n289_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT27), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n280_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n276_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n299_), .A2(KEYINPUT20), .A3(new_n267_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(KEYINPUT97), .A2(new_n298_), .B1(new_n300_), .B2(new_n294_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n253_), .A2(new_n266_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n290_), .A2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n303_), .B(KEYINPUT20), .C1(new_n290_), .C2(new_n276_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT97), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n280_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n288_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT98), .B1(new_n297_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n288_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT20), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n310_), .B1(new_n290_), .B2(new_n276_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n294_), .B1(new_n311_), .B2(new_n267_), .ZN(new_n312_));
  OAI22_X1  g111(.A1(new_n312_), .A2(KEYINPUT94), .B1(new_n304_), .B2(new_n280_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n289_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n296_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  AND2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT1), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT85), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(G141gat), .B2(G148gat), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .A4(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n325_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n327_), .B(KEYINPUT3), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n329_), .B(KEYINPUT2), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n324_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n321_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n319_), .B(new_n320_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n324_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n327_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n329_), .B(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n339_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n338_), .B(new_n344_), .C1(new_n325_), .C2(new_n332_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n337_), .A2(new_n345_), .A3(KEYINPUT4), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT95), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n321_), .B(new_n349_), .C1(new_n333_), .C2(new_n336_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n337_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n352_));
  INV_X1    g151(.A(G85gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT0), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G57gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(G57gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n353_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n355_), .A2(G57gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(G85gat), .A3(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n351_), .A2(new_n352_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n298_), .A2(KEYINPUT97), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n300_), .A2(new_n294_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n306_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n309_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT98), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT27), .A4(new_n296_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n308_), .A2(new_n318_), .A3(new_n365_), .A4(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT29), .B1(new_n333_), .B2(new_n336_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n290_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT87), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(G228gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(G228gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n290_), .A2(new_n382_), .A3(new_n373_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G78gat), .B(G106gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT93), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n333_), .A2(new_n336_), .A3(KEYINPUT29), .ZN(new_n388_));
  XOR2_X1   g187(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n389_));
  XNOR2_X1  g188(.A(G22gat), .B(G50gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n388_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n385_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n381_), .A2(new_n383_), .A3(new_n393_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n387_), .A2(new_n392_), .B1(new_n394_), .B2(new_n386_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n396_));
  AND4_X1   g195(.A1(new_n396_), .A2(new_n386_), .A3(new_n394_), .A4(new_n392_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G15gat), .B(G43gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT83), .Z(new_n401_));
  INV_X1    g200(.A(KEYINPUT30), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n245_), .A2(new_n252_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n258_), .A2(new_n265_), .A3(new_n241_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n266_), .B(KEYINPUT30), .C1(new_n245_), .C2(new_n252_), .ZN(new_n406_));
  INV_X1    g205(.A(G227gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n375_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n405_), .A2(new_n406_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n401_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT30), .B1(new_n253_), .B2(new_n266_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n406_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n408_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n405_), .A2(new_n406_), .A3(new_n409_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n401_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G71gat), .B(G99gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n412_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n419_), .B1(new_n412_), .B2(new_n418_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT31), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n412_), .A2(new_n418_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n419_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT31), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n427_), .A2(new_n421_), .A3(new_n428_), .A4(new_n420_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n424_), .A2(new_n321_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n321_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n399_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n424_), .A2(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n338_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n424_), .A2(new_n321_), .A3(new_n429_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n398_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n372_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n288_), .A2(KEYINPUT32), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n365_), .B1(new_n368_), .B2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n283_), .A2(new_n438_), .A3(new_n289_), .A4(new_n295_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT96), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n281_), .A2(new_n282_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT96), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n438_), .A4(new_n289_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n346_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n337_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(new_n361_), .A3(new_n359_), .A4(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n363_), .B2(KEYINPUT33), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n351_), .A2(new_n352_), .A3(new_n362_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n296_), .A3(new_n315_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n446_), .A2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n456_), .B(new_n398_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n437_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G57gat), .B(G64gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n460_), .A2(KEYINPUT11), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(KEYINPUT11), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G71gat), .B(G78gat), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(new_n463_), .A3(KEYINPUT11), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT68), .ZN(new_n467_));
  XOR2_X1   g266(.A(G15gat), .B(G22gat), .Z(new_n468_));
  NAND2_X1  g267(.A1(G1gat), .A2(G8gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(KEYINPUT14), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT73), .ZN(new_n471_));
  XOR2_X1   g270(.A(G1gat), .B(G8gat), .Z(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n470_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n472_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(KEYINPUT74), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(KEYINPUT74), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G231gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(new_n375_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n481_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n486_), .A2(new_n483_), .A3(new_n375_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n467_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G183gat), .B(G211gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(G127gat), .B(G155gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n493_), .A2(KEYINPUT17), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n482_), .A2(new_n484_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n486_), .B1(new_n483_), .B2(new_n375_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n467_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n488_), .A2(new_n494_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n488_), .A2(KEYINPUT76), .A3(new_n494_), .A4(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n485_), .A2(new_n487_), .A3(new_n466_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n466_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n493_), .A2(KEYINPUT17), .ZN(new_n507_));
  OR4_X1    g306(.A1(new_n504_), .A2(new_n506_), .A3(new_n494_), .A4(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G85gat), .B(G92gat), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n515_));
  NOR2_X1   g314(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n516_));
  OAI22_X1  g315(.A1(new_n515_), .A2(new_n516_), .B1(G99gat), .B2(G106gat), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n514_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(KEYINPUT66), .A3(new_n520_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n511_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n521_), .A2(new_n514_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n510_), .A2(new_n526_), .ZN(new_n528_));
  OAI22_X1  g327(.A1(new_n525_), .A2(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G29gat), .B(G36gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G43gat), .B(G50gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n353_), .A2(new_n287_), .A3(KEYINPUT9), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n514_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT10), .B(G99gat), .Z(new_n536_));
  INV_X1    g335(.A(KEYINPUT64), .ZN(new_n537_));
  INV_X1    g336(.A(G106gat), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n533_), .B(new_n535_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n529_), .A2(new_n532_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT65), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT7), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n518_), .B1(new_n545_), .B2(new_n519_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n518_), .A2(new_n519_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n522_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n514_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n524_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n526_), .B1(new_n550_), .B2(new_n510_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n527_), .A2(new_n528_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n541_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n532_), .B(KEYINPUT15), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT71), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT34), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT35), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n542_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(new_n559_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT36), .ZN(new_n567_));
  INV_X1    g366(.A(new_n562_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n542_), .A2(new_n555_), .A3(new_n568_), .A4(new_n560_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n563_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT72), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n563_), .A2(new_n569_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n566_), .B(KEYINPUT36), .Z(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT37), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n459_), .A2(new_n509_), .A3(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n466_), .B(new_n541_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT67), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n553_), .A2(new_n505_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n467_), .A2(KEYINPUT12), .A3(new_n553_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n581_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n586_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT69), .B1(new_n584_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT69), .ZN(new_n593_));
  AOI211_X1 g392(.A(new_n593_), .B(KEYINPUT12), .C1(new_n553_), .C2(new_n505_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n588_), .B(new_n590_), .C1(new_n592_), .C2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n212_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT5), .B(G176gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  NAND3_X1  g398(.A1(new_n587_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT70), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n587_), .A2(new_n595_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n599_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n602_), .B(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT13), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n605_), .B1(new_n601_), .B2(new_n600_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n608_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n473_), .A2(new_n477_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n532_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n532_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n478_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G229gat), .A2(G233gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n618_), .B(KEYINPUT77), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n478_), .A2(new_n554_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n614_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(G169gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n211_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n620_), .A2(new_n624_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n620_), .B2(new_n624_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT78), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n620_), .A2(new_n624_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n627_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT78), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(new_n628_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT79), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT79), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n580_), .A2(new_n612_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(G1gat), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n365_), .B(KEYINPUT99), .Z(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n644_), .A2(new_n645_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT38), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT100), .B1(new_n612_), .B2(new_n637_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n652_), .B(new_n638_), .C1(new_n607_), .C2(new_n611_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n509_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n575_), .B(KEYINPUT101), .Z(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n459_), .ZN(new_n658_));
  AND4_X1   g457(.A1(new_n651_), .A2(new_n654_), .A3(new_n655_), .A4(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n365_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n649_), .B1(new_n645_), .B2(new_n661_), .ZN(G1324gat));
  INV_X1    g461(.A(G8gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n308_), .A2(new_n318_), .A3(new_n371_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n659_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(KEYINPUT39), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(KEYINPUT39), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n644_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT103), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n668_), .A2(new_n674_), .A3(new_n670_), .A4(new_n671_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n673_), .A2(KEYINPUT40), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT40), .B1(new_n673_), .B2(new_n675_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n430_), .A2(new_n431_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n659_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT41), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n644_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1326gat));
  INV_X1    g483(.A(G22gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n659_), .B2(new_n399_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT104), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT42), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n644_), .A2(new_n685_), .A3(new_n399_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n459_), .A2(new_n656_), .ZN(new_n691_));
  AND4_X1   g490(.A1(new_n612_), .A2(new_n691_), .A3(new_n509_), .A4(new_n642_), .ZN(new_n692_));
  INV_X1    g491(.A(G29gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n660_), .A2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT106), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n579_), .B1(new_n437_), .B2(new_n458_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(KEYINPUT43), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(KEYINPUT43), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n579_), .B(new_n702_), .C1(new_n437_), .C2(new_n458_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n700_), .A2(new_n701_), .A3(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n651_), .A2(new_n654_), .A3(new_n509_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n697_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n701_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n698_), .A2(new_n699_), .A3(KEYINPUT43), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n703_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n650_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(KEYINPUT44), .A3(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n707_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(new_n647_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n696_), .B1(new_n714_), .B2(new_n693_), .ZN(G1328gat));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n664_), .A3(new_n712_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n707_), .A2(new_n712_), .A3(KEYINPUT107), .A4(new_n664_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(G36gat), .A3(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(G36gat), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n664_), .A2(KEYINPUT108), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n664_), .A2(KEYINPUT108), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n692_), .A2(new_n721_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n720_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n720_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n730_), .A2(KEYINPUT46), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n721_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT109), .B(new_n727_), .C1(new_n735_), .C2(new_n719_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n731_), .B1(new_n720_), .B2(new_n728_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n733_), .A2(new_n738_), .ZN(G1329gat));
  AOI21_X1  g538(.A(G43gat), .B1(new_n692_), .B2(new_n680_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n680_), .A2(G43gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n713_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g542(.A(G50gat), .B1(new_n692_), .B2(new_n399_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n399_), .A2(G50gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n713_), .B2(new_n745_), .ZN(G1331gat));
  NOR2_X1   g545(.A1(new_n612_), .A2(new_n637_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n580_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n646_), .B1(new_n748_), .B2(KEYINPUT110), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(KEYINPUT110), .B2(new_n748_), .ZN(new_n750_));
  INV_X1    g549(.A(G57gat), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n639_), .A2(new_n503_), .A3(new_n508_), .A4(new_n641_), .ZN(new_n752_));
  NOR4_X1   g551(.A1(new_n657_), .A2(new_n752_), .A3(new_n459_), .A4(new_n612_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n365_), .A2(new_n751_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n750_), .A2(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1332gat));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n753_), .B2(new_n724_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT48), .Z(new_n758_));
  INV_X1    g557(.A(new_n748_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(new_n756_), .A3(new_n724_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1333gat));
  INV_X1    g560(.A(G71gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n753_), .B2(new_n680_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT49), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n762_), .A3(new_n680_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT111), .Z(G1334gat));
  INV_X1    g566(.A(G78gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n753_), .B2(new_n399_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT50), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n759_), .A2(new_n768_), .A3(new_n399_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1335gat));
  OR2_X1    g571(.A1(new_n710_), .A2(KEYINPUT112), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n710_), .A2(KEYINPUT112), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n655_), .A2(new_n612_), .A3(new_n637_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n365_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n775_), .A2(new_n691_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n353_), .A3(new_n647_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1336gat));
  INV_X1    g579(.A(new_n724_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G92gat), .B1(new_n776_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(new_n287_), .A3(new_n664_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1337gat));
  INV_X1    g583(.A(new_n680_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G99gat), .B1(new_n776_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n778_), .A2(new_n536_), .A3(new_n680_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT51), .ZN(G1338gat));
  AND2_X1   g588(.A1(new_n775_), .A2(new_n399_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n538_), .B1(new_n710_), .B2(new_n790_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT52), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n538_), .A3(new_n691_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g594(.A1(new_n752_), .A2(new_n579_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n612_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n796_), .B2(new_n612_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n614_), .A2(new_n623_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n622_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n803_), .B2(new_n802_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n627_), .B1(new_n617_), .B2(new_n622_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n629_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n606_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n637_), .A2(new_n600_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n583_), .B(new_n588_), .C1(new_n592_), .C2(new_n594_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n586_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n595_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n466_), .B1(new_n529_), .B2(new_n541_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n593_), .B1(new_n814_), .B2(KEYINPUT12), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n584_), .A2(KEYINPUT69), .A3(new_n591_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(KEYINPUT55), .A3(new_n588_), .A4(new_n590_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n811_), .A2(new_n813_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n811_), .A2(new_n813_), .A3(new_n818_), .A4(KEYINPUT114), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n604_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n599_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT56), .A3(new_n822_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n809_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n808_), .B1(new_n828_), .B2(KEYINPUT115), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n830_), .B(new_n809_), .C1(new_n825_), .C2(new_n827_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n656_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT57), .B(new_n656_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n579_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n825_), .A2(new_n837_), .A3(new_n827_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n807_), .A2(new_n600_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n826_), .B2(new_n822_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(KEYINPUT117), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n836_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n838_), .A2(new_n841_), .A3(KEYINPUT58), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n834_), .A2(new_n835_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n801_), .B1(new_n847_), .B2(new_n509_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n436_), .A2(new_n664_), .A3(new_n646_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n637_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT59), .B1(new_n848_), .B2(new_n850_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n832_), .A2(new_n833_), .B1(new_n845_), .B2(new_n844_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n655_), .B1(new_n856_), .B2(new_n835_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n855_), .B(new_n849_), .C1(new_n857_), .C2(new_n801_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n854_), .A2(new_n858_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n859_), .A2(new_n642_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n853_), .B1(new_n860_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g660(.A(new_n612_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n854_), .A2(new_n862_), .A3(new_n858_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G120gat), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865_));
  AOI21_X1  g664(.A(G120gat), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n865_), .B2(G120gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n851_), .A2(KEYINPUT118), .A3(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n849_), .B(new_n867_), .C1(new_n857_), .C2(new_n801_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n864_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT119), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n864_), .A2(new_n875_), .A3(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1341gat));
  INV_X1    g676(.A(G127gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n851_), .A2(new_n878_), .A3(new_n655_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n859_), .A2(new_n655_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n878_), .ZN(G1342gat));
  AOI21_X1  g680(.A(G134gat), .B1(new_n851_), .B2(new_n657_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n882_), .A2(KEYINPUT120), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(KEYINPUT120), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n579_), .A2(G134gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT121), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n883_), .A2(new_n884_), .B1(new_n859_), .B2(new_n886_), .ZN(G1343gat));
  NOR2_X1   g686(.A1(new_n848_), .A2(new_n432_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(new_n647_), .A3(new_n781_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n638_), .ZN(new_n890_));
  INV_X1    g689(.A(G141gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n612_), .ZN(new_n893_));
  INV_X1    g692(.A(G148gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1345gat));
  NOR2_X1   g694(.A1(new_n889_), .A2(new_n509_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT61), .B(G155gat), .Z(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  NAND2_X1  g697(.A1(new_n579_), .A2(G162gat), .ZN(new_n899_));
  XOR2_X1   g698(.A(new_n899_), .B(KEYINPUT123), .Z(new_n900_));
  NOR2_X1   g699(.A1(new_n889_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(G162gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n889_), .B2(new_n656_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT122), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n905_), .B(new_n902_), .C1(new_n889_), .C2(new_n656_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n901_), .B1(new_n904_), .B2(new_n906_), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n848_), .A2(new_n399_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n724_), .A2(new_n680_), .A3(new_n646_), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(KEYINPUT124), .Z(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911_), .B2(new_n638_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT62), .B(G169gat), .C1(new_n911_), .C2(new_n638_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n911_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n916_), .A2(new_n637_), .A3(new_n272_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n915_), .A3(new_n917_), .ZN(G1348gat));
  OR2_X1    g717(.A1(new_n908_), .A2(KEYINPUT125), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n908_), .A2(KEYINPUT125), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n862_), .A2(G176gat), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n919_), .A2(new_n910_), .A3(new_n920_), .A4(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n271_), .B1(new_n911_), .B2(new_n612_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1349gat));
  NAND4_X1  g723(.A1(new_n919_), .A2(new_n655_), .A3(new_n910_), .A4(new_n920_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n509_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n925_), .A2(new_n230_), .B1(new_n916_), .B2(new_n926_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n911_), .B2(new_n836_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n657_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n911_), .B2(new_n929_), .ZN(G1351gat));
  NOR2_X1   g729(.A1(new_n781_), .A2(new_n660_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n888_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n638_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n211_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n612_), .ZN(new_n935_));
  MUX2_X1   g734(.A(G204gat), .B(new_n214_), .S(new_n935_), .Z(G1353gat));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n205_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n655_), .B1(new_n937_), .B2(new_n205_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT126), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n888_), .A2(new_n931_), .A3(new_n938_), .A4(new_n941_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n937_), .B(new_n205_), .C1(new_n932_), .C2(new_n940_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n942_), .A2(KEYINPUT127), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(G1354gat));
  OAI21_X1  g745(.A(G218gat), .B1(new_n932_), .B2(new_n836_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n657_), .A2(new_n207_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n932_), .B2(new_n948_), .ZN(G1355gat));
endmodule


