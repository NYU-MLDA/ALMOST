//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT85), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n204_), .A2(KEYINPUT85), .A3(G183gat), .A4(G190gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(G169gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT26), .B(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n217_), .A2(KEYINPUT24), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n203_), .A2(new_n205_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n213_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G120gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(G127gat), .A2(G134gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G127gat), .A2(G134gat), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n226_), .A2(new_n227_), .A3(G113gat), .ZN(new_n228_));
  INV_X1    g027(.A(G113gat), .ZN(new_n229_));
  INV_X1    g028(.A(G127gat), .ZN(new_n230_));
  INV_X1    g029(.A(G134gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G127gat), .A2(G134gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n229_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n225_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(G113gat), .B1(new_n226_), .B2(new_n227_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(G120gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n224_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G15gat), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT31), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n240_), .B(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G99gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  XNOR2_X1  g046(.A(new_n243_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n250_));
  OR2_X1    g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT87), .B1(new_n254_), .B2(KEYINPUT86), .ZN(new_n255_));
  OR2_X1    g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n257_));
  OAI22_X1  g056(.A1(new_n255_), .A2(new_n256_), .B1(new_n257_), .B2(KEYINPUT3), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT86), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n257_), .B1(new_n262_), .B2(KEYINPUT3), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n261_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n258_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT88), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n253_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n252_), .A2(KEYINPUT1), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(G155gat), .A3(G162gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n273_), .A3(new_n251_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G141gat), .B(G148gat), .Z(new_n275_));
  AND2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n239_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n255_), .A2(new_n256_), .B1(new_n260_), .B2(new_n259_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n257_), .A2(KEYINPUT3), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n269_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n253_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n276_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n236_), .A2(new_n237_), .A3(G120gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(G120gat), .B1(new_n236_), .B2(new_n237_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT96), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT96), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n235_), .A2(new_n287_), .A3(new_n238_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n250_), .B1(new_n277_), .B2(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n284_), .A2(new_n285_), .A3(KEYINPUT96), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT97), .B1(new_n293_), .B2(new_n283_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n290_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT98), .B(G85gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G29gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT0), .B(G57gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n239_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(new_n283_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(KEYINPUT4), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n283_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT97), .B1(new_n308_), .B2(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n289_), .A2(new_n250_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n307_), .B1(new_n311_), .B2(KEYINPUT4), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n298_), .B(new_n304_), .C1(new_n312_), .C2(new_n295_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT4), .B1(new_n290_), .B2(new_n294_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n307_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n295_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n303_), .B1(new_n316_), .B2(new_n297_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G233gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT89), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(G228gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(G228gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n319_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n283_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT90), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(G204gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(KEYINPUT21), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G197gat), .B(G204gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n334_), .A2(KEYINPUT21), .A3(new_n327_), .A4(new_n330_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n327_), .A2(KEYINPUT21), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n324_), .B1(new_n326_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n324_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n339_), .B(new_n340_), .C1(new_n283_), .C2(new_n325_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G78gat), .B(G106gat), .Z(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n338_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n283_), .A2(new_n325_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT28), .B(G22gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G50gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n348_), .B(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n343_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(KEYINPUT91), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n345_), .A2(KEYINPUT91), .A3(new_n346_), .A4(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT19), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT92), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n221_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT94), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n220_), .A2(KEYINPUT93), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT94), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n221_), .A2(new_n207_), .A3(new_n364_), .A4(new_n209_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n216_), .A2(new_n366_), .A3(new_n219_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n222_), .A2(new_n208_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n212_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n337_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT20), .B1(new_n339_), .B2(new_n224_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n360_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT18), .ZN(new_n375_));
  INV_X1    g174(.A(G64gat), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n376_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n377_), .A2(G92gat), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(G92gat), .B1(new_n377_), .B2(new_n378_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n368_), .A2(new_n337_), .A3(new_n370_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n339_), .B2(new_n224_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n384_), .A3(new_n359_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n373_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n381_), .B1(new_n373_), .B2(new_n385_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n357_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n381_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n371_), .A2(new_n372_), .A3(new_n360_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n359_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n373_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(KEYINPUT27), .A3(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n318_), .A2(KEYINPUT100), .A3(new_n356_), .A4(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT100), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n356_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n313_), .A2(new_n317_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT99), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(KEYINPUT33), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n313_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n314_), .A2(new_n315_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n297_), .B1(new_n405_), .B2(new_n296_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n403_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n304_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n295_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n409_), .B(new_n303_), .C1(new_n295_), .C2(new_n311_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n373_), .A2(new_n385_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n389_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(KEYINPUT95), .A3(new_n393_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n404_), .A2(new_n408_), .A3(new_n410_), .A4(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n390_), .A2(new_n391_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n419_), .A2(new_n413_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n399_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n356_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n249_), .B1(new_n401_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT101), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT101), .B(new_n249_), .C1(new_n401_), .C2(new_n423_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n249_), .A2(new_n399_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n395_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n429_), .A2(new_n356_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n426_), .A2(new_n427_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G230gat), .A2(G233gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT68), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G99gat), .ZN(new_n438_));
  INV_X1    g237(.A(G106gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT6), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(G99gat), .A3(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT68), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n434_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n437_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G85gat), .ZN(new_n449_));
  INV_X1    g248(.A(G92gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G85gat), .A2(G92gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT67), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n448_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n448_), .A2(KEYINPUT69), .A3(new_n457_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(KEYINPUT8), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n443_), .A2(new_n434_), .A3(new_n445_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n457_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n450_), .A2(KEYINPUT64), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT64), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G92gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n469_), .A3(G85gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n451_), .A2(KEYINPUT9), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT65), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT10), .B(G99gat), .Z(new_n480_));
  AOI22_X1  g279(.A1(new_n480_), .A2(new_n439_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n479_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G71gat), .B(G78gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G71gat), .B(G78gat), .Z(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(KEYINPUT11), .A3(new_n486_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT70), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n466_), .A2(new_n485_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n484_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n433_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT71), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n493_), .B(KEYINPUT72), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT12), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n495_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT73), .B(KEYINPUT12), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n496_), .B2(new_n494_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n432_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT71), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(new_n433_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n499_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G120gat), .B(G148gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT5), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(G176gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(G204gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT74), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n499_), .A2(new_n506_), .A3(new_n513_), .A4(new_n508_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522_));
  INV_X1    g321(.A(G169gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(new_n329_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G29gat), .B(G36gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G43gat), .A2(G50gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G43gat), .A2(G50gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT77), .B1(new_n536_), .B2(new_n531_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n530_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n530_), .B1(new_n537_), .B2(new_n535_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n528_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n529_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n530_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n527_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT83), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n540_), .A2(new_n544_), .A3(KEYINPUT83), .ZN(new_n548_));
  INV_X1    g347(.A(G15gat), .ZN(new_n549_));
  INV_X1    g348(.A(G22gat), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(G15gat), .A2(G22gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(G1gat), .A2(G8gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT14), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT80), .B1(new_n553_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT80), .ZN(new_n558_));
  OAI221_X1 g357(.A(new_n558_), .B1(new_n554_), .B2(new_n555_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(G1gat), .A2(G8gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n554_), .A2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n557_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n547_), .A2(new_n548_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT84), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n547_), .A2(KEYINPUT84), .A3(new_n548_), .A4(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n547_), .A2(new_n548_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n526_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n526_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n540_), .A2(new_n544_), .A3(KEYINPUT15), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT15), .B1(new_n540_), .B2(new_n544_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n564_), .ZN(new_n577_));
  AOI211_X1 g376(.A(new_n574_), .B(new_n577_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n525_), .B1(new_n573_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n569_), .A2(new_n526_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n525_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n567_), .A2(new_n568_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n581_), .B(new_n582_), .C1(new_n526_), .C2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n521_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n431_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n466_), .A2(new_n545_), .A3(new_n485_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n576_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n540_), .A2(new_n544_), .A3(KEYINPUT15), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n591_), .B(new_n596_), .C1(new_n599_), .C2(new_n496_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT79), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n496_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n591_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n594_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n496_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n575_), .A2(new_n576_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT79), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n591_), .A4(new_n596_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n601_), .A2(new_n604_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT78), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(G134gat), .ZN(new_n613_));
  INV_X1    g412(.A(G162gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n610_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n610_), .B2(new_n618_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n590_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n601_), .A2(new_n609_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n622_), .A2(new_n616_), .A3(new_n615_), .A4(new_n604_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n610_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(KEYINPUT37), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n564_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n564_), .A2(new_n627_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(new_n494_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G127gat), .B(G155gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT17), .Z(new_n637_));
  NOR2_X1   g436(.A1(new_n631_), .A2(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n630_), .A2(new_n500_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n630_), .A2(new_n500_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n639_), .A2(KEYINPUT17), .A3(new_n640_), .A4(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT82), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n643_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n638_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n626_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n589_), .A2(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n649_), .A2(G1gat), .A3(new_n318_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(KEYINPUT103), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT103), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n652_), .B(new_n653_), .Z(new_n654_));
  NOR2_X1   g453(.A1(new_n619_), .A2(new_n620_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n431_), .A2(KEYINPUT104), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT104), .B1(new_n431_), .B2(new_n655_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n656_), .A2(new_n587_), .A3(new_n646_), .A4(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n318_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(G1324gat));
  OR3_X1    g459(.A1(new_n649_), .A2(G8gat), .A3(new_n395_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n656_), .A2(new_n646_), .A3(new_n657_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(new_n587_), .A3(new_n429_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(G8gat), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n662_), .B(G8gat), .C1(new_n658_), .C2(new_n395_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n661_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT40), .B(new_n661_), .C1(new_n665_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(new_n649_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n549_), .A3(new_n248_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G15gat), .B1(new_n658_), .B2(new_n249_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT105), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(KEYINPUT105), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(KEYINPUT41), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n676_), .B2(new_n677_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n674_), .B1(new_n678_), .B2(new_n679_), .ZN(G1326gat));
  NAND3_X1  g479(.A1(new_n673_), .A2(new_n550_), .A3(new_n356_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n663_), .A2(new_n587_), .A3(new_n356_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(G22gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n682_), .B2(G22gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n681_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  NOR3_X1   g486(.A1(new_n646_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n589_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G29gat), .B1(new_n689_), .B2(new_n399_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n587_), .A2(new_n647_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n430_), .A2(new_n428_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n407_), .B1(new_n406_), .B2(new_n304_), .ZN(new_n695_));
  NOR4_X1   g494(.A1(new_n316_), .A2(new_n297_), .A3(new_n303_), .A4(new_n403_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n311_), .A2(new_n295_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n295_), .B2(new_n405_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n303_), .A2(new_n699_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n313_), .A2(new_n317_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n701_));
  AOI22_X1  g500(.A1(new_n697_), .A2(new_n700_), .B1(new_n701_), .B2(new_n421_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n400_), .B(new_n396_), .C1(new_n702_), .C2(new_n356_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT101), .B1(new_n703_), .B2(new_n249_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n427_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n694_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n626_), .B(KEYINPUT106), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n693_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n626_), .A2(new_n693_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n431_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n692_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT44), .B(new_n692_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n399_), .A2(G29gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n690_), .B1(new_n716_), .B2(new_n717_), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n714_), .A2(new_n429_), .A3(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT107), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n714_), .A2(new_n721_), .A3(new_n429_), .A4(new_n715_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(G36gat), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724_));
  INV_X1    g523(.A(G36gat), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n689_), .A2(new_n724_), .A3(new_n725_), .A4(new_n429_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n589_), .A2(new_n725_), .A3(new_n688_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT108), .B1(new_n727_), .B2(new_n395_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n726_), .A2(KEYINPUT45), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT45), .B1(new_n726_), .B2(new_n728_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n723_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n723_), .A2(new_n733_), .A3(new_n731_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1329gat));
  NAND2_X1  g536(.A1(new_n689_), .A2(new_n248_), .ZN(new_n738_));
  XOR2_X1   g537(.A(KEYINPUT111), .B(G43gat), .Z(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n714_), .A2(G43gat), .A3(new_n248_), .A4(new_n715_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT110), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT110), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT47), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(new_n740_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1330gat));
  INV_X1    g547(.A(G50gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n689_), .A2(new_n749_), .A3(new_n356_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n716_), .A2(new_n356_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n749_), .ZN(G1331gat));
  OR2_X1    g551(.A1(new_n519_), .A2(new_n520_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(new_n585_), .ZN(new_n754_));
  AND4_X1   g553(.A1(G57gat), .A2(new_n663_), .A3(new_n399_), .A4(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n431_), .A2(new_n585_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT112), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(new_n521_), .A3(new_n648_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n399_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(G57gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n755_), .B1(new_n762_), .B2(new_n763_), .ZN(G1332gat));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n376_), .A3(new_n429_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n663_), .A2(new_n429_), .A3(new_n754_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(G64gat), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n766_), .B2(G64gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n765_), .B1(new_n769_), .B2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n758_), .A2(new_n772_), .A3(new_n248_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n663_), .A2(new_n248_), .A3(new_n754_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(G71gat), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n774_), .B2(G71gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(new_n777_), .B2(new_n778_), .ZN(G1334gat));
  INV_X1    g578(.A(G78gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n758_), .A2(new_n780_), .A3(new_n356_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n663_), .A2(new_n356_), .A3(new_n754_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(G78gat), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n782_), .B2(G78gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n781_), .B1(new_n785_), .B2(new_n786_), .ZN(G1335gat));
  NAND2_X1  g586(.A1(new_n754_), .A2(new_n647_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT114), .Z(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT43), .B1(new_n431_), .B2(new_n707_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n706_), .A2(new_n693_), .A3(new_n626_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n792_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n793_), .A2(new_n449_), .A3(new_n318_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n757_), .A2(new_n521_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(new_n688_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n399_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n794_), .B1(new_n797_), .B2(new_n449_), .ZN(G1336gat));
  AOI21_X1  g597(.A(G92gat), .B1(new_n796_), .B2(new_n429_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n793_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n429_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(G1337gat));
  AND2_X1   g601(.A1(new_n248_), .A2(new_n480_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n795_), .A2(new_n688_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n438_), .B1(new_n800_), .B2(new_n248_), .ZN(new_n805_));
  OR3_X1    g604(.A1(new_n804_), .A2(KEYINPUT51), .A3(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT51), .B1(new_n804_), .B2(new_n805_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1338gat));
  INV_X1    g607(.A(new_n356_), .ZN(new_n809_));
  OAI21_X1  g608(.A(G106gat), .B1(new_n793_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT115), .B(G106gat), .C1(new_n793_), .C2(new_n809_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(KEYINPUT52), .A3(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n795_), .A2(new_n439_), .A3(new_n356_), .A4(new_n688_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n810_), .A2(new_n811_), .A3(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT53), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n814_), .A2(new_n820_), .A3(new_n815_), .A4(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1339gat));
  NAND2_X1  g621(.A1(new_n585_), .A2(new_n518_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT117), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n585_), .A2(new_n825_), .A3(new_n518_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n432_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n506_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n503_), .A2(KEYINPUT55), .A3(new_n432_), .A4(new_n505_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n831_), .B2(new_n515_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n833_), .B(new_n514_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n824_), .B(new_n826_), .C1(new_n832_), .C2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n516_), .A2(new_n518_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n569_), .A2(new_n574_), .A3(new_n580_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n837_), .B(new_n525_), .C1(new_n574_), .C2(new_n583_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n838_), .A2(new_n584_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n655_), .B1(new_n835_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT57), .B1(new_n841_), .B2(KEYINPUT118), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n518_), .B(new_n839_), .C1(new_n832_), .C2(new_n834_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n621_), .A2(new_n625_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n518_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n496_), .A2(new_n501_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n496_), .A2(new_n494_), .ZN(new_n851_));
  AND4_X1   g650(.A1(new_n432_), .A2(new_n850_), .A3(new_n851_), .A4(new_n505_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n851_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n505_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n433_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n852_), .B1(new_n855_), .B2(KEYINPUT55), .ZN(new_n856_));
  INV_X1    g655(.A(new_n830_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n515_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n833_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n831_), .A2(KEYINPUT56), .A3(new_n515_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n849_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n861_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n839_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n846_), .A2(new_n848_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n585_), .A2(new_n825_), .A3(new_n518_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n825_), .B1(new_n585_), .B2(new_n518_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n859_), .A2(new_n860_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n868_), .A2(new_n869_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n864_), .B(new_n865_), .C1(new_n870_), .C2(new_n655_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n842_), .A2(new_n863_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n647_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n621_), .A2(new_n625_), .A3(new_n586_), .A4(new_n646_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n874_), .A2(new_n521_), .A3(KEYINPUT116), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT116), .B1(new_n874_), .B2(new_n521_), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT54), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n877_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n879_), .A2(new_n875_), .A3(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n873_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n429_), .A2(new_n318_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n248_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n883_), .A2(new_n809_), .A3(new_n885_), .A4(new_n888_), .ZN(new_n889_));
  AOI211_X1 g688(.A(new_n356_), .B(new_n887_), .C1(new_n873_), .C2(new_n882_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n885_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n889_), .B1(new_n890_), .B2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n586_), .A2(new_n229_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(KEYINPUT121), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G113gat), .B1(new_n896_), .B2(KEYINPUT121), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n585_), .A3(new_n890_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1340gat));
  AOI21_X1  g698(.A(new_n356_), .B1(new_n873_), .B2(new_n882_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n225_), .A2(KEYINPUT60), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n225_), .B1(new_n753_), .B2(KEYINPUT60), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n900_), .A2(new_n888_), .A3(new_n901_), .A4(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n890_), .A2(KEYINPUT122), .A3(new_n901_), .A4(new_n902_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n225_), .B1(new_n894_), .B2(new_n521_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT123), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n906_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n883_), .A2(new_n809_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n892_), .B1(new_n912_), .B2(new_n887_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n753_), .B1(new_n913_), .B2(new_n889_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n910_), .B(new_n911_), .C1(new_n914_), .C2(new_n225_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n909_), .A2(new_n915_), .ZN(G1341gat));
  AOI21_X1  g715(.A(G127gat), .B1(new_n890_), .B2(new_n646_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n647_), .B1(new_n913_), .B2(new_n889_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g718(.A(G134gat), .B1(new_n890_), .B2(new_n655_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT124), .B(G134gat), .Z(new_n921_));
  NOR2_X1   g720(.A1(new_n847_), .A2(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n894_), .B2(new_n922_), .ZN(G1343gat));
  AOI211_X1 g722(.A(new_n248_), .B(new_n809_), .C1(new_n873_), .C2(new_n882_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n924_), .A2(new_n886_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n585_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n521_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n646_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT61), .B(G155gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1346gat));
  AOI21_X1  g731(.A(G162gat), .B1(new_n925_), .B2(new_n655_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n707_), .A2(new_n614_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n925_), .B2(new_n934_), .ZN(G1347gat));
  NAND4_X1  g734(.A1(new_n900_), .A2(new_n585_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n937_));
  OAI21_X1  g736(.A(G169gat), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n936_), .B2(KEYINPUT22), .ZN(new_n939_));
  MUX2_X1   g738(.A(G169gat), .B(new_n938_), .S(new_n939_), .Z(G1348gat));
  AND3_X1   g739(.A1(new_n900_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n521_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT126), .B(G176gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1349gat));
  NAND2_X1  g743(.A1(new_n941_), .A2(new_n646_), .ZN(new_n945_));
  MUX2_X1   g744(.A(new_n214_), .B(G183gat), .S(new_n945_), .Z(G1350gat));
  NAND3_X1  g745(.A1(new_n941_), .A2(new_n655_), .A3(new_n215_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n941_), .A2(new_n626_), .ZN(new_n948_));
  INV_X1    g747(.A(G190gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n947_), .B1(new_n948_), .B2(new_n949_), .ZN(G1351gat));
  NOR2_X1   g749(.A1(new_n395_), .A2(new_n399_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n924_), .A2(new_n951_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n952_), .A2(new_n586_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(new_n329_), .ZN(G1352gat));
  INV_X1    g753(.A(new_n952_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n521_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  AND2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  NOR4_X1   g758(.A1(new_n952_), .A2(new_n647_), .A3(new_n958_), .A4(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n955_), .A2(new_n646_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n961_), .B2(new_n958_), .ZN(G1354gat));
  AOI21_X1  g761(.A(G218gat), .B1(new_n955_), .B2(new_n655_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n626_), .A2(G218gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(KEYINPUT127), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n955_), .B2(new_n965_), .ZN(G1355gat));
endmodule


