//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  AOI22_X1  g002(.A1(new_n202_), .A2(new_n203_), .B1(G71gat), .B2(G78gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT69), .B1(new_n202_), .B2(new_n203_), .ZN(new_n205_));
  INV_X1    g004(.A(G71gat), .ZN(new_n206_));
  INV_X1    g005(.A(G78gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G57gat), .B(G64gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT11), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n205_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n208_), .B(new_n213_), .C1(new_n209_), .C2(KEYINPUT11), .ZN(new_n214_));
  INV_X1    g013(.A(new_n211_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n210_), .B1(new_n209_), .B2(KEYINPUT11), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(G231gat), .A2(G233gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G8gat), .ZN(new_n222_));
  INV_X1    g021(.A(G1gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT79), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT79), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G1gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n226_), .A3(G8gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT14), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n229_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n232_), .A2(G1gat), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n230_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT80), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n223_), .B1(new_n236_), .B2(new_n231_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n222_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(G1gat), .B1(new_n232_), .B2(new_n233_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n223_), .A3(new_n231_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(G8gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n221_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G127gat), .B(G155gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT16), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G183gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(G211gat), .Z(new_n247_));
  INV_X1    g046(.A(KEYINPUT17), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n243_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n243_), .A2(new_n249_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G232gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT34), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n255_), .A2(KEYINPUT35), .ZN(new_n256_));
  XOR2_X1   g055(.A(G29gat), .B(G36gat), .Z(new_n257_));
  INV_X1    g056(.A(KEYINPUT75), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G29gat), .B(G36gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT75), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G43gat), .ZN(new_n263_));
  INV_X1    g062(.A(G43gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n264_), .A3(new_n261_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n263_), .A2(G50gat), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(G50gat), .B1(new_n263_), .B2(new_n265_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT10), .B(G99gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n270_));
  OR3_X1    g069(.A1(new_n269_), .A2(new_n270_), .A3(G106gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(G85gat), .B(G92gat), .Z(new_n272_));
  NAND2_X1  g071(.A1(G99gat), .A2(G106gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT6), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(G99gat), .A3(G106gat), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n272_), .A2(KEYINPUT9), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G85gat), .ZN(new_n278_));
  INV_X1    g077(.A(G92gat), .ZN(new_n279_));
  OR3_X1    g078(.A1(new_n278_), .A2(new_n279_), .A3(KEYINPUT9), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n270_), .B1(new_n269_), .B2(G106gat), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n271_), .A2(new_n277_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT7), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G99gat), .A2(G106gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n274_), .A2(new_n276_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n286_), .A2(KEYINPUT67), .A3(new_n287_), .A4(new_n288_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .A4(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n272_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT8), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT8), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n299_), .A2(new_n304_), .A3(new_n301_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n283_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT76), .B(KEYINPUT15), .Z(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT77), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n299_), .A2(new_n304_), .A3(new_n301_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n304_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n282_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n268_), .B1(new_n308_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n307_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n268_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n256_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n306_), .A2(KEYINPUT77), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n317_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n308_), .A2(new_n268_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n255_), .A2(KEYINPUT35), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n256_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n319_), .A2(new_n320_), .A3(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G190gat), .B(G218gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G134gat), .ZN(new_n329_));
  INV_X1    g128(.A(G162gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT36), .ZN(new_n333_));
  INV_X1    g132(.A(new_n331_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n319_), .A2(new_n326_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n327_), .A2(KEYINPUT36), .A3(new_n331_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT37), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(KEYINPUT37), .A3(new_n337_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(KEYINPUT22), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G169gat), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n344_), .B(new_n347_), .C1(new_n348_), .C2(new_n345_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353_));
  MUX2_X1   g152(.A(new_n352_), .B(KEYINPUT23), .S(new_n353_), .Z(new_n354_));
  NOR2_X1   g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n349_), .A2(new_n350_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n351_), .A2(new_n357_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT25), .B(G183gat), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n367_), .B2(new_n358_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n352_), .B1(G183gat), .B2(G190gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n353_), .A2(KEYINPUT23), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n364_), .B(new_n368_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n360_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT86), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT86), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n360_), .A2(new_n374_), .A3(new_n371_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT31), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT30), .Z(new_n378_));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379_));
  INV_X1    g178(.A(G113gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G120gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(new_n206_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n382_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G15gat), .B(G43gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT87), .B(G99gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n378_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT105), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n394_), .B(new_n395_), .Z(new_n396_));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n397_), .B(KEYINPUT92), .Z(new_n398_));
  XOR2_X1   g197(.A(new_n398_), .B(KEYINPUT19), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G197gat), .B(G204gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT21), .ZN(new_n404_));
  XOR2_X1   g203(.A(G211gat), .B(G218gat), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT21), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n402_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n401_), .B2(KEYINPUT91), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n410_), .B(new_n405_), .C1(KEYINPUT91), .C2(new_n401_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n356_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n348_), .A2(new_n344_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n358_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT93), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n363_), .B(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n368_), .B(new_n354_), .C1(new_n417_), .C2(new_n361_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n412_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n376_), .B2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n400_), .B1(new_n422_), .B2(KEYINPUT20), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n415_), .A2(new_n418_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n425_), .A2(KEYINPUT20), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n376_), .B2(new_n421_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n427_), .A2(new_n399_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n396_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n360_), .A2(new_n374_), .A3(new_n371_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n374_), .B1(new_n360_), .B2(new_n371_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n421_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(KEYINPUT20), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n399_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n396_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n421_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n419_), .A2(KEYINPUT94), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n412_), .A2(new_n415_), .A3(new_n438_), .A4(new_n418_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n436_), .A2(KEYINPUT20), .A3(new_n440_), .A4(new_n400_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n434_), .A2(new_n435_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT103), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT103), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n434_), .A2(new_n441_), .A3(new_n444_), .A4(new_n435_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n429_), .A2(new_n443_), .A3(KEYINPUT27), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT104), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n436_), .A2(KEYINPUT20), .A3(new_n419_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n399_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n427_), .B2(new_n399_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n449_), .B1(new_n452_), .B2(new_n396_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n453_), .A2(KEYINPUT104), .A3(new_n443_), .A4(new_n445_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n434_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n441_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n396_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT27), .B1(new_n458_), .B2(new_n442_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n382_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G155gat), .A2(G162gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G155gat), .A2(G162gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G141gat), .A2(G148gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT2), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n463_), .B(new_n464_), .C1(new_n467_), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n465_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n464_), .B(KEYINPUT1), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n472_), .B(new_n468_), .C1(new_n473_), .C2(new_n462_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n471_), .A2(KEYINPUT96), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n461_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(KEYINPUT88), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n382_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n471_), .A2(new_n474_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(KEYINPUT88), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n476_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n482_), .A2(KEYINPUT100), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n479_), .B(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT97), .B(KEYINPUT4), .Z(new_n488_));
  OR3_X1    g287(.A1(new_n487_), .A2(new_n461_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT4), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n489_), .B(new_n484_), .C1(new_n482_), .C2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT100), .B1(new_n482_), .B2(new_n484_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n485_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT99), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G29gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G85gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n485_), .A2(new_n491_), .A3(new_n501_), .A4(new_n492_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G228gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT89), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT29), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n421_), .B(new_n505_), .C1(new_n487_), .C2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n412_), .B1(KEYINPUT29), .B2(new_n479_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G22gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n509_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n487_), .A2(new_n506_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G50gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n516_), .B(G50gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n512_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n503_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  AND4_X1   g321(.A1(new_n391_), .A2(new_n455_), .A3(new_n460_), .A4(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n459_), .B1(new_n448_), .B2(new_n454_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n391_), .B1(new_n524_), .B2(new_n522_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n502_), .A2(KEYINPUT33), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n502_), .A2(KEYINPUT33), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n442_), .B(new_n458_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n499_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT101), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n489_), .B(new_n483_), .C1(new_n490_), .C2(new_n482_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT102), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n452_), .A2(KEYINPUT32), .A3(new_n435_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n503_), .A2(new_n537_), .ZN(new_n538_));
  AOI211_X1 g337(.A(new_n457_), .B(new_n456_), .C1(KEYINPUT32), .C2(new_n435_), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n529_), .A2(new_n536_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n519_), .A2(new_n521_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n390_), .B1(new_n526_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n503_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n524_), .A2(new_n390_), .A3(new_n545_), .A4(new_n542_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n253_), .B(new_n343_), .C1(new_n544_), .C2(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n238_), .A2(new_n268_), .A3(new_n241_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n268_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n315_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n317_), .A2(new_n307_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT81), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT81), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n558_), .B(new_n555_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT82), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n346_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(G197gat), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n554_), .A2(new_n557_), .A3(new_n559_), .A4(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n282_), .B(new_n218_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT12), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n303_), .A2(new_n305_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n218_), .B1(new_n573_), .B2(new_n282_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n576_));
  INV_X1    g375(.A(new_n218_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n311_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n570_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n570_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n571_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n587_), .B1(new_n574_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n311_), .A2(new_n577_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n571_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT70), .A3(new_n587_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n580_), .A2(new_n586_), .A3(new_n591_), .A4(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(KEYINPUT12), .A3(new_n571_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n587_), .B1(new_n596_), .B2(new_n578_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT70), .B1(new_n593_), .B2(new_n587_), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n590_), .B(new_n570_), .C1(new_n592_), .C2(new_n571_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n585_), .B(KEYINPUT72), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n595_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT73), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n580_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT73), .B1(new_n605_), .B2(new_n601_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT13), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n606_), .B1(new_n603_), .B2(KEYINPUT73), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT13), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT74), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n548_), .A2(new_n569_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n224_), .A2(new_n226_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n503_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n455_), .A2(new_n460_), .A3(new_n522_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT105), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n524_), .A2(new_n391_), .A3(new_n522_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n543_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n390_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n547_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n613_), .A2(new_n568_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n336_), .A2(KEYINPUT106), .A3(new_n337_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT106), .B1(new_n336_), .B2(new_n337_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n253_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n545_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n618_), .A2(new_n619_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n620_), .A2(new_n635_), .A3(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT107), .ZN(new_n639_));
  INV_X1    g438(.A(new_n524_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n628_), .A2(new_n640_), .A3(new_n633_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G8gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT39), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n644_), .A3(G8gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n524_), .A2(G8gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n615_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n639_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n641_), .A2(new_n644_), .A3(G8gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n644_), .B1(new_n641_), .B2(G8gat), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n648_), .B(new_n639_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n638_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n648_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT107), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(KEYINPUT40), .A3(new_n652_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(G1325gat));
  INV_X1    g457(.A(G15gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n615_), .A2(new_n659_), .A3(new_n390_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n628_), .A2(new_n390_), .A3(new_n633_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n661_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(new_n661_), .B2(G15gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n660_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT108), .Z(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n615_), .A2(new_n666_), .A3(new_n541_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n634_), .B2(new_n542_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT109), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT109), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(KEYINPUT42), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT42), .B1(new_n669_), .B2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(new_n671_), .B2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n338_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n336_), .A2(KEYINPUT106), .A3(new_n337_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n253_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n628_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G29gat), .B1(new_n679_), .B2(new_n503_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n681_), .B(new_n342_), .C1(new_n544_), .C2(new_n547_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT43), .B1(new_n626_), .B2(new_n343_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n627_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n685_), .A4(new_n632_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n686_), .A2(G29gat), .A3(new_n503_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n685_), .A3(new_n632_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n680_), .B1(new_n687_), .B2(new_n690_), .ZN(G1328gat));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  AOI211_X1 g492(.A(new_n627_), .B(new_n253_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n524_), .B1(new_n694_), .B2(KEYINPUT44), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n695_), .B2(new_n690_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n679_), .A2(new_n693_), .A3(new_n640_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n692_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n694_), .A2(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n686_), .A2(new_n640_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G36gat), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(KEYINPUT46), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n705_), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n690_), .A2(G43gat), .A3(new_n390_), .A4(new_n686_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n679_), .A2(new_n390_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n264_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT47), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1330gat));
  NAND3_X1  g513(.A1(new_n690_), .A2(new_n541_), .A3(new_n686_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G50gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n541_), .A2(new_n517_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT110), .Z(new_n718_));
  NAND2_X1  g517(.A1(new_n679_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1331gat));
  NOR2_X1   g519(.A1(new_n613_), .A2(new_n568_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n548_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n503_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n614_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n626_), .A2(new_n568_), .A3(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n633_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(KEYINPUT111), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(KEYINPUT111), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n503_), .A2(G57gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n724_), .B1(new_n730_), .B2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n723_), .A2(new_n733_), .A3(new_n640_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n728_), .A2(new_n640_), .A3(new_n729_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G64gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G64gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n723_), .A2(new_n206_), .A3(new_n390_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n728_), .A2(new_n390_), .A3(new_n729_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT49), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G71gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G71gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1334gat));
  NAND3_X1  g544(.A1(new_n723_), .A2(new_n207_), .A3(new_n541_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n728_), .A2(new_n541_), .A3(new_n729_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(G78gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G78gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n726_), .A2(new_n678_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n503_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n253_), .B(new_n722_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n545_), .A2(new_n278_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  OAI21_X1  g556(.A(new_n279_), .B1(new_n752_), .B2(new_n524_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n758_), .A2(KEYINPUT112), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(KEYINPUT112), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(G92gat), .A3(new_n640_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT113), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n759_), .A2(new_n764_), .A3(new_n760_), .A4(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1337gat));
  NAND2_X1  g565(.A1(new_n755_), .A2(new_n390_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G99gat), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n752_), .A2(new_n269_), .A3(new_n625_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT51), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n768_), .A2(new_n769_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1338gat));
  OR3_X1    g573(.A1(new_n752_), .A2(G106gat), .A3(new_n542_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n684_), .A2(new_n541_), .A3(new_n632_), .A4(new_n721_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G106gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n775_), .B(new_n782_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1339gat));
  NOR2_X1   g583(.A1(new_n608_), .A2(KEYINPUT13), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n610_), .A2(new_n611_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n341_), .B(new_n340_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n253_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT114), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT54), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n788_), .B(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n343_), .A2(new_n791_), .A3(new_n613_), .A4(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n790_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n596_), .A2(new_n578_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n570_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n580_), .A2(KEYINPUT55), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n597_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n797_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n602_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n597_), .A2(new_n799_), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT55), .B(new_n587_), .C1(new_n596_), .C2(new_n578_), .ZN(new_n805_));
  OAI22_X1  g604(.A1(new_n804_), .A2(new_n805_), .B1(new_n570_), .B2(new_n796_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT56), .B1(new_n806_), .B2(new_n601_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n568_), .B(new_n595_), .C1(new_n803_), .C2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n551_), .A2(new_n555_), .A3(new_n553_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n552_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n565_), .A3(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n567_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n608_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n808_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n677_), .A2(new_n814_), .A3(KEYINPUT57), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n802_), .B1(new_n801_), .B2(new_n602_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n601_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n567_), .A2(new_n595_), .A3(new_n811_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(KEYINPUT58), .A3(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n342_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n815_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n566_), .A2(new_n567_), .B1(new_n586_), .B2(new_n600_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n818_), .A2(new_n827_), .B1(new_n608_), .B2(new_n812_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n631_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT115), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n826_), .C1(new_n631_), .C2(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n825_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n795_), .B1(new_n833_), .B2(new_n632_), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n640_), .A2(new_n625_), .A3(new_n545_), .A4(new_n541_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837_), .B2(new_n568_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n829_), .A2(new_n815_), .A3(new_n824_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n632_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n840_), .B2(new_n632_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n795_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n839_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT59), .B1(new_n834_), .B2(new_n836_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n840_), .A2(new_n632_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT116), .ZN(new_n850_));
  INV_X1    g649(.A(new_n795_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n840_), .A2(new_n841_), .A3(new_n632_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(KEYINPUT117), .A3(new_n845_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n847_), .A2(new_n848_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n569_), .A2(new_n380_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n838_), .B1(new_n855_), .B2(new_n856_), .ZN(G1340gat));
  NAND4_X1  g656(.A1(new_n847_), .A2(new_n614_), .A3(new_n848_), .A4(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G120gat), .ZN(new_n859_));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n613_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n837_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n860_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT118), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n859_), .A2(new_n865_), .A3(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1341gat));
  AOI21_X1  g666(.A(G127gat), .B1(new_n837_), .B2(new_n253_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n253_), .A2(G127gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n855_), .B2(new_n869_), .ZN(G1342gat));
  XOR2_X1   g669(.A(KEYINPUT119), .B(G134gat), .Z(new_n871_));
  NOR2_X1   g670(.A1(new_n343_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n847_), .A2(new_n848_), .A3(new_n854_), .A4(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n834_), .A2(new_n677_), .A3(new_n836_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(G134gat), .B2(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT120), .ZN(G1343gat));
  NOR3_X1   g675(.A1(new_n834_), .A2(new_n390_), .A3(new_n542_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n640_), .A2(new_n545_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n877_), .A2(KEYINPUT121), .A3(new_n878_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n568_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G141gat), .ZN(new_n885_));
  INV_X1    g684(.A(G141gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n886_), .A3(new_n568_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n883_), .A2(new_n614_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G148gat), .ZN(new_n890_));
  INV_X1    g689(.A(G148gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n883_), .A2(new_n891_), .A3(new_n614_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n883_), .A2(new_n253_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT122), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n883_), .A2(new_n253_), .A3(new_n896_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1346gat));
  AOI21_X1  g699(.A(G162gat), .B1(new_n883_), .B2(new_n631_), .ZN(new_n901_));
  AOI211_X1 g700(.A(new_n330_), .B(new_n343_), .C1(new_n881_), .C2(new_n882_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1347gat));
  NOR4_X1   g702(.A1(new_n625_), .A2(new_n524_), .A3(new_n503_), .A4(new_n541_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n853_), .A2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905_), .B2(new_n569_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT123), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n906_), .A2(new_n909_), .A3(KEYINPUT62), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n905_), .B(KEYINPUT124), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n568_), .A2(new_n348_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT125), .ZN(new_n915_));
  OAI22_X1  g714(.A1(new_n911_), .A2(new_n912_), .B1(new_n913_), .B2(new_n915_), .ZN(G1348gat));
  OR2_X1    g715(.A1(new_n913_), .A2(new_n613_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n834_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(new_n904_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n725_), .A2(new_n344_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n917_), .A2(new_n344_), .B1(new_n919_), .B2(new_n920_), .ZN(G1349gat));
  NOR3_X1   g720(.A1(new_n913_), .A2(new_n362_), .A3(new_n632_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G183gat), .B1(new_n919_), .B2(new_n253_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n913_), .B2(new_n343_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n677_), .A2(new_n417_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n913_), .B2(new_n926_), .ZN(G1351gat));
  NOR2_X1   g726(.A1(new_n834_), .A2(new_n390_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n928_), .A2(new_n640_), .A3(new_n522_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n568_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n614_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G204gat), .ZN(G1353gat));
  OAI22_X1  g733(.A1(new_n929_), .A2(new_n632_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  XOR2_X1   g735(.A(KEYINPUT63), .B(G211gat), .Z(new_n937_));
  NOR3_X1   g736(.A1(new_n929_), .A2(new_n632_), .A3(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(KEYINPUT126), .B1(new_n936_), .B2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n930_), .A2(new_n253_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n935_), .B(new_n940_), .C1(new_n941_), .C2(new_n937_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n939_), .A2(new_n942_), .ZN(G1354gat));
  OR3_X1    g742(.A1(new_n929_), .A2(KEYINPUT127), .A3(new_n677_), .ZN(new_n944_));
  INV_X1    g743(.A(G218gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(KEYINPUT127), .B1(new_n929_), .B2(new_n677_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n944_), .A2(new_n945_), .A3(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n930_), .A2(G218gat), .A3(new_n342_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1355gat));
endmodule


