//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n215_), .B2(KEYINPUT2), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT3), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n214_), .A2(KEYINPUT91), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n216_), .A2(new_n219_), .A3(new_n221_), .A4(new_n222_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT90), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n212_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n212_), .B(KEYINPUT92), .C1(new_n225_), .C2(new_n223_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n209_), .B1(KEYINPUT1), .B2(new_n210_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n210_), .A2(KEYINPUT1), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n232_), .B(KEYINPUT89), .Z(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n215_), .A2(new_n217_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n206_), .B1(new_n237_), .B2(KEYINPUT99), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n228_), .A2(new_n229_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT99), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n205_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n202_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT100), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n202_), .A3(new_n205_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  OR3_X1    g046(.A1(new_n242_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n243_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n238_), .A2(new_n241_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n245_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n248_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G1gat), .B(G29gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G57gat), .B(G85gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n249_), .A2(new_n251_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n257_), .A3(new_n248_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G8gat), .B(G36gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT22), .B(G169gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n276_), .B2(G176gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT82), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281_));
  MUX2_X1   g080(.A(new_n278_), .B(new_n280_), .S(new_n281_), .Z(new_n282_));
  NOR2_X1   g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n277_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(KEYINPUT24), .A3(new_n274_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT25), .B(G183gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n281_), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT84), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(new_n281_), .B2(new_n280_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n288_), .A2(KEYINPUT24), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT97), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n293_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT97), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n285_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G197gat), .B(G204gat), .Z(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(KEYINPUT21), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(KEYINPUT21), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n273_), .B1(new_n302_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT102), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n282_), .A2(new_n297_), .A3(new_n292_), .A4(new_n289_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n296_), .A2(new_n284_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n275_), .A2(KEYINPUT83), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT83), .B1(new_n316_), .B2(G169gat), .ZN(new_n317_));
  INV_X1    g116(.A(G176gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n274_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n313_), .B1(new_n314_), .B2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n311_), .A2(new_n312_), .B1(new_n309_), .B2(new_n321_), .ZN(new_n322_));
  AOI211_X1 g121(.A(new_n309_), .B(new_n285_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT102), .B1(new_n323_), .B2(new_n273_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n272_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n296_), .B2(new_n284_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n297_), .A2(new_n292_), .A3(new_n289_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(new_n282_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n273_), .B1(new_n328_), .B2(new_n310_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n310_), .B2(new_n302_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(new_n271_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n269_), .B1(new_n325_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT103), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT103), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(new_n269_), .C1(new_n325_), .C2(new_n331_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n271_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n271_), .B1(new_n321_), .B2(new_n309_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n311_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n339_), .A3(new_n268_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n262_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT33), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n261_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n260_), .A2(KEYINPUT33), .A3(new_n257_), .A4(new_n248_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n267_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n300_), .A2(new_n301_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n309_), .B1(new_n346_), .B2(new_n285_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n272_), .B1(new_n347_), .B2(new_n329_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n321_), .A2(new_n309_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n272_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n350_), .A2(new_n323_), .A3(new_n273_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n345_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n337_), .A2(new_n339_), .A3(new_n267_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n244_), .A2(new_n245_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n242_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n257_), .B1(new_n250_), .B2(new_n246_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n343_), .A2(new_n344_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n310_), .B1(new_n237_), .B2(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G228gat), .A2(G233gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT93), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n361_), .A2(KEYINPUT93), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  OAI221_X1 g165(.A(new_n309_), .B1(new_n363_), .B2(new_n365_), .C1(new_n239_), .C2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G78gat), .B(G106gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT94), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G22gat), .B(G50gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n239_), .B2(new_n366_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n239_), .A2(new_n374_), .A3(new_n366_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n373_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n377_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n373_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n380_), .A2(new_n375_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n364_), .A2(new_n367_), .A3(new_n370_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n372_), .A2(new_n384_), .A3(KEYINPUT95), .A4(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT95), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n378_), .A2(new_n382_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n367_), .B(new_n391_), .C1(new_n360_), .C2(new_n363_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n389_), .B(new_n369_), .C1(new_n392_), .C2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n386_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n341_), .A2(new_n359_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n398_), .B(G15gat), .Z(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT85), .B(G43gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n328_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n321_), .A2(new_n404_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n401_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n205_), .B(KEYINPUT31), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n328_), .A2(new_n405_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n321_), .A2(new_n404_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n400_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n413_), .A2(KEYINPUT86), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(KEYINPUT86), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n409_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT87), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI211_X1 g217(.A(KEYINPUT87), .B(new_n409_), .C1(new_n408_), .C2(new_n412_), .ZN(new_n419_));
  OAI22_X1  g218(.A1(new_n414_), .A2(new_n415_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT27), .B1(new_n352_), .B2(new_n353_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n345_), .B1(new_n325_), .B2(new_n331_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n353_), .A2(KEYINPUT27), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n261_), .A3(new_n259_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n396_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n420_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n396_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n259_), .A2(new_n261_), .A3(new_n420_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT104), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n259_), .A2(new_n261_), .A3(new_n420_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT104), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n396_), .A4(new_n424_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n397_), .A2(new_n427_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G29gat), .B(G36gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G43gat), .B(G50gat), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G43gat), .B(G50gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT14), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT74), .B(G8gat), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(G1gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(G15gat), .B(G22gat), .Z(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT75), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(KEYINPUT74), .A2(G8gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(KEYINPUT74), .A2(G8gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(G1gat), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT14), .ZN(new_n450_));
  INV_X1    g249(.A(new_n445_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G1gat), .B(G8gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n446_), .B2(new_n453_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n441_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n446_), .A2(new_n453_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT68), .B(KEYINPUT15), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n438_), .A2(new_n440_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n465_), .A3(new_n455_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT79), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n461_), .A2(new_n455_), .A3(new_n440_), .A4(new_n438_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n458_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT79), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n458_), .A2(new_n466_), .A3(new_n474_), .A4(new_n467_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G113gat), .B(G141gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G169gat), .B(G197gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  NAND4_X1  g277(.A1(new_n469_), .A2(new_n473_), .A3(new_n475_), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT80), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n468_), .A2(KEYINPUT79), .B1(new_n471_), .B2(new_n472_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n475_), .A4(new_n478_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n475_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n478_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n434_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  AND4_X1   g298(.A1(new_n493_), .A2(new_n497_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT66), .ZN(new_n501_));
  AND2_X1   g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G85gat), .ZN(new_n505_));
  INV_X1    g304(.A(G92gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G85gat), .A2(G92gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT66), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT8), .B1(new_n500_), .B2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n497_), .A2(new_n493_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT8), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n504_), .A4(new_n509_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n516_));
  OR2_X1    g315(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(KEYINPUT64), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT64), .ZN(new_n520_));
  AND2_X1   g319(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n496_), .ZN(new_n525_));
  AND3_X1   g324(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n507_), .A2(KEYINPUT9), .A3(new_n508_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n508_), .A2(KEYINPUT9), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n516_), .B1(new_n525_), .B2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(G106gat), .B1(new_n519_), .B2(new_n523_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n533_), .A2(new_n534_), .A3(KEYINPUT65), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n515_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT67), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n539_));
  XOR2_X1   g338(.A(G71gat), .B(G78gat), .Z(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n525_), .A2(new_n531_), .A3(new_n516_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT65), .B1(new_n533_), .B2(new_n534_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT67), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n515_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n537_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n544_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n536_), .A2(KEYINPUT12), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n544_), .B1(new_n537_), .B2(new_n549_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n550_), .B(new_n552_), .C1(new_n553_), .C2(KEYINPUT12), .ZN(new_n554_));
  AND2_X1   g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n549_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n548_), .B1(new_n547_), .B2(new_n515_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n551_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n550_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n555_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n557_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n557_), .B2(new_n562_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT13), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n461_), .A2(new_n455_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n461_), .B2(new_n455_), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n544_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n544_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n579_), .B1(new_n585_), .B2(KEYINPUT76), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(KEYINPUT76), .B2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT77), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT77), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n586_), .B(new_n589_), .C1(KEYINPUT76), .C2(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n585_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n576_), .B(KEYINPUT17), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT78), .B1(new_n591_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT78), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n598_), .B(new_n595_), .C1(new_n588_), .C2(new_n590_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT71), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT36), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT72), .Z(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n537_), .A2(new_n441_), .A3(new_n549_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT70), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n537_), .A2(KEYINPUT70), .A3(new_n441_), .A4(new_n549_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n536_), .A2(new_n465_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT69), .Z(new_n617_));
  AOI21_X1  g416(.A(new_n610_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n610_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n607_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n615_), .A2(new_n617_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n610_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n621_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n605_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n622_), .A2(KEYINPUT73), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT73), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n607_), .B(new_n629_), .C1(new_n618_), .C2(new_n621_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT37), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n625_), .A2(new_n627_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n632_), .A2(KEYINPUT37), .A3(new_n622_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n572_), .A2(new_n601_), .A3(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n490_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(G1gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n262_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n622_), .A2(KEYINPUT73), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n642_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n434_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n591_), .A2(new_n596_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n572_), .A2(new_n489_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n262_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n639_), .A2(new_n640_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n641_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT105), .Z(G1324gat));
  INV_X1    g451(.A(new_n637_), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n653_), .A2(new_n424_), .A3(new_n443_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G8gat), .B1(new_n647_), .B2(new_n424_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(KEYINPUT39), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(KEYINPUT39), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n654_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n658_), .B(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(new_n420_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G15gat), .B1(new_n647_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n653_), .A2(G15gat), .A3(new_n662_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  OAI21_X1  g465(.A(G22gat), .B1(new_n647_), .B2(new_n396_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT42), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n396_), .A2(G22gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n653_), .B2(new_n669_), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n601_), .A2(new_n643_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n572_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n490_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G29gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n262_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n572_), .A2(new_n489_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n601_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n434_), .B2(new_n634_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n397_), .A2(new_n427_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n430_), .A2(new_n433_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n635_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n677_), .B1(new_n678_), .B2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n262_), .B1(new_n684_), .B2(KEYINPUT44), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n682_), .B1(new_n681_), .B2(new_n635_), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT43), .B(new_n634_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n601_), .B(new_n676_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n684_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n685_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G29gat), .B1(new_n693_), .B2(new_n694_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n675_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n424_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n673_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT45), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n684_), .A2(KEYINPUT44), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n424_), .B(new_n703_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT46), .B(new_n702_), .C1(new_n704_), .C2(new_n699_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n691_), .A2(new_n692_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n703_), .A2(new_n424_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n699_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n701_), .B(KEYINPUT45), .Z(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n705_), .A2(new_n711_), .ZN(G1329gat));
  AOI21_X1  g511(.A(G43gat), .B1(new_n673_), .B2(new_n420_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n691_), .A2(new_n692_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n703_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(G43gat), .A3(new_n420_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n714_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT47), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(new_n714_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1330gat));
  AOI21_X1  g521(.A(G50gat), .B1(new_n673_), .B2(new_n426_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n716_), .A2(G50gat), .A3(new_n426_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n707_), .ZN(G1331gat));
  NOR3_X1   g524(.A1(new_n601_), .A2(new_n571_), .A3(new_n488_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n644_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(G57gat), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n648_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n434_), .A2(new_n488_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n601_), .A2(new_n635_), .A3(new_n571_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n648_), .B1(new_n733_), .B2(KEYINPUT109), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(KEYINPUT109), .B2(new_n733_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n729_), .B1(new_n735_), .B2(new_n728_), .ZN(G1332gat));
  OAI21_X1  g535(.A(G64gat), .B1(new_n727_), .B2(new_n424_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT48), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n424_), .A2(G64gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n732_), .B2(new_n739_), .ZN(G1333gat));
  OR3_X1    g539(.A1(new_n732_), .A2(G71gat), .A3(new_n662_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n644_), .A2(new_n420_), .A3(new_n726_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G71gat), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n743_), .A2(KEYINPUT111), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(KEYINPUT111), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n741_), .B1(new_n747_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n727_), .B2(new_n396_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n396_), .A2(G78gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n732_), .B2(new_n752_), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n671_), .A2(new_n571_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n730_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n505_), .A3(new_n262_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n678_), .A2(new_n683_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n571_), .A2(new_n600_), .A3(new_n488_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n262_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n761_), .B2(new_n505_), .ZN(G1336gat));
  NAND3_X1  g561(.A1(new_n756_), .A2(new_n506_), .A3(new_n700_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n760_), .A2(new_n700_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n506_), .ZN(G1337gat));
  AND3_X1   g564(.A1(new_n756_), .A2(new_n420_), .A3(new_n524_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n760_), .A2(new_n420_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G99gat), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g568(.A1(new_n756_), .A2(new_n496_), .A3(new_n426_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n426_), .B(new_n759_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n758_), .A2(KEYINPUT112), .A3(new_n426_), .A4(new_n759_), .ZN(new_n774_));
  XOR2_X1   g573(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n775_));
  AND4_X1   g574(.A1(G106gat), .A2(new_n773_), .A3(new_n774_), .A4(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n496_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n777_), .B2(new_n774_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n770_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n770_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  NOR2_X1   g582(.A1(new_n648_), .A2(new_n662_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n428_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n645_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n556_), .B1(new_n555_), .B2(new_n561_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n791_), .A2(new_n567_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n555_), .A2(KEYINPUT114), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n554_), .B2(new_n793_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n550_), .A2(new_n552_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT12), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n560_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n798_), .A2(new_n800_), .A3(KEYINPUT55), .A4(new_n795_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n797_), .A3(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n566_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n792_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n471_), .A2(new_n467_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n458_), .A2(new_n466_), .A3(new_n472_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n486_), .A3(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n484_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n643_), .B1(new_n805_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n789_), .B(new_n790_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n628_), .A2(new_n630_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n557_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n488_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n802_), .A2(new_n566_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n810_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n814_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT117), .B1(new_n823_), .B2(KEYINPUT115), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT57), .B1(new_n811_), .B2(new_n789_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n813_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n815_), .A2(new_n484_), .A3(new_n808_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n828_), .A2(KEYINPUT58), .B1(new_n631_), .B2(new_n633_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n829_), .A2(new_n830_), .B1(KEYINPUT58), .B2(new_n828_), .ZN(new_n831_));
  OAI221_X1 g630(.A(KEYINPUT116), .B1(new_n631_), .B2(new_n633_), .C1(KEYINPUT58), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n788_), .B1(new_n826_), .B2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n571_), .A2(new_n600_), .A3(new_n489_), .A4(new_n634_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n787_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G113gat), .B1(new_n839_), .B2(new_n488_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n790_), .B1(new_n823_), .B2(KEYINPUT117), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n789_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n844_), .A2(new_n813_), .B1(new_n832_), .B2(new_n831_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n845_), .B2(new_n600_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n835_), .B(KEYINPUT54), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n826_), .A2(new_n833_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(KEYINPUT120), .A3(new_n601_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n786_), .B2(KEYINPUT119), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(KEYINPUT119), .B2(new_n786_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT121), .B1(new_n850_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n600_), .B1(new_n826_), .B2(new_n833_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n847_), .B1(new_n856_), .B2(KEYINPUT120), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n845_), .A2(new_n841_), .A3(new_n600_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT121), .B(new_n853_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT118), .B1(new_n838_), .B2(KEYINPUT59), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n838_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n855_), .A2(new_n859_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n488_), .A2(G113gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n840_), .B1(new_n863_), .B2(new_n864_), .ZN(G1340gat));
  INV_X1    g664(.A(new_n859_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n854_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n838_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n572_), .B1(new_n868_), .B2(new_n860_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G120gat), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n571_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n839_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n871_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n839_), .B2(new_n600_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n788_), .A2(G127gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n863_), .B2(new_n876_), .ZN(G1342gat));
  AOI21_X1  g676(.A(G134gat), .B1(new_n839_), .B2(new_n643_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n635_), .A2(G134gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n863_), .B2(new_n879_), .ZN(G1343gat));
  OAI21_X1  g679(.A(new_n847_), .B1(new_n845_), .B2(new_n788_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n396_), .A2(new_n420_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n648_), .A2(new_n700_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n489_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT122), .B(G141gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1344gat));
  NOR2_X1   g686(.A1(new_n884_), .A2(new_n571_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g688(.A1(new_n884_), .A2(new_n601_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT61), .B(G155gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  OR3_X1    g691(.A1(new_n884_), .A2(G162gat), .A3(new_n814_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G162gat), .B1(new_n884_), .B2(new_n634_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n893_), .A2(new_n894_), .A3(KEYINPUT123), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n262_), .A2(new_n424_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n420_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n426_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n850_), .A2(new_n488_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G169gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n905_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n903_), .A2(new_n276_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(G1348gat));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n850_), .A2(new_n572_), .A3(new_n902_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n912_), .B2(G176gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(KEYINPUT125), .A3(new_n318_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n881_), .A2(new_n396_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n571_), .A2(new_n901_), .A3(new_n318_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n913_), .A2(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1349gat));
  NOR2_X1   g716(.A1(new_n601_), .A2(new_n901_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n915_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(G183gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n645_), .A2(new_n290_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n850_), .A2(new_n902_), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT126), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n921_), .A2(new_n926_), .A3(new_n923_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n850_), .A2(new_n635_), .A3(new_n902_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G190gat), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n850_), .A2(new_n291_), .A3(new_n643_), .A4(new_n902_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(KEYINPUT127), .A3(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1351gat));
  AND2_X1   g735(.A1(new_n881_), .A2(new_n882_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n937_), .A2(new_n488_), .A3(new_n900_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g738(.A1(new_n937_), .A2(new_n572_), .A3(new_n900_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g740(.A(KEYINPUT63), .B(G211gat), .ZN(new_n942_));
  OR2_X1    g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n937_), .A2(new_n788_), .A3(new_n900_), .ZN(new_n944_));
  MUX2_X1   g743(.A(new_n942_), .B(new_n943_), .S(new_n944_), .Z(G1354gat));
  NAND2_X1  g744(.A1(new_n937_), .A2(new_n900_), .ZN(new_n946_));
  OAI21_X1  g745(.A(G218gat), .B1(new_n946_), .B2(new_n634_), .ZN(new_n947_));
  OR2_X1    g746(.A1(new_n814_), .A2(G218gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n946_), .B2(new_n948_), .ZN(G1355gat));
endmodule


