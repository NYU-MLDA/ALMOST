//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n968_, new_n969_, new_n971_, new_n972_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n999_, new_n1000_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n207_));
  OAI22_X1  g006(.A1(new_n206_), .A2(new_n207_), .B1(G85gat), .B2(G92gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(new_n207_), .B2(new_n206_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT65), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT10), .B(G99gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n216_), .B(new_n217_), .C1(new_n218_), .C2(G106gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT66), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT67), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n221_), .A2(new_n223_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT68), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n223_), .A4(new_n221_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n216_), .A2(new_n217_), .A3(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT69), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G85gat), .B(G92gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT70), .B(KEYINPUT8), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n236_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT8), .B1(new_n237_), .B2(new_n240_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n220_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G29gat), .B(G36gat), .Z(new_n246_));
  XOR2_X1   g045(.A(G43gat), .B(G50gat), .Z(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G232gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT35), .Z(new_n254_));
  OAI21_X1  g053(.A(new_n242_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n255_));
  AOI211_X1 g054(.A(KEYINPUT69), .B(new_n235_), .C1(new_n229_), .C2(new_n232_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n244_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT73), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT73), .B(new_n244_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n220_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n248_), .B(KEYINPUT15), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n250_), .B(new_n254_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n220_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(new_n248_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT73), .B1(new_n243_), .B2(new_n244_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n260_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n264_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n262_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n266_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n253_), .A2(KEYINPUT35), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n205_), .B(new_n263_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT76), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n250_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT35), .A3(new_n253_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n205_), .A4(new_n263_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n263_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n204_), .B(KEYINPUT36), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n279_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G15gat), .B(G22gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT78), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n289_), .A2(new_n290_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n290_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT79), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G15gat), .B(G22gat), .Z(new_n298_));
  INV_X1    g097(.A(KEYINPUT14), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(G1gat), .B2(G8gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT78), .B1(new_n298_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(new_n294_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G1gat), .B(G8gat), .Z(new_n304_));
  NAND3_X1  g103(.A1(new_n297_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n297_), .B2(new_n303_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(G231gat), .A2(G233gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n308_), .A2(new_n309_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(KEYINPUT71), .A2(G71gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(KEYINPUT71), .A2(G71gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G78gat), .ZN(new_n317_));
  INV_X1    g116(.A(G78gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n318_), .A3(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT11), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G57gat), .B(G64gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(KEYINPUT11), .A3(new_n319_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n323_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n317_), .A2(KEYINPUT11), .A3(new_n319_), .A4(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n313_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n313_), .A2(new_n330_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G127gat), .B(G155gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(G183gat), .B(G211gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n337_), .A2(KEYINPUT17), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n332_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT81), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n325_), .A2(new_n328_), .A3(KEYINPUT72), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT72), .B1(new_n325_), .B2(new_n328_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n311_), .A2(new_n344_), .A3(new_n312_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n337_), .A2(KEYINPUT17), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n345_), .A2(new_n338_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n343_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n325_), .A2(new_n328_), .A3(KEYINPUT72), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n350_), .B2(new_n313_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n339_), .A2(new_n340_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n341_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n288_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G57gat), .B(G85gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT103), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G1gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n358_));
  INV_X1    g157(.A(G29gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n357_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  OR2_X1    g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n362_), .B1(new_n363_), .B2(KEYINPUT3), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT2), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(G141gat), .A3(G148gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(KEYINPUT3), .ZN(new_n370_));
  NOR2_X1   g169(.A1(G141gat), .A2(G148gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(KEYINPUT90), .A3(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n364_), .A2(new_n369_), .A3(new_n370_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(KEYINPUT1), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(G155gat), .A3(G162gat), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n378_), .A2(new_n380_), .A3(new_n376_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT89), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n371_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n365_), .A3(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n377_), .A2(KEYINPUT91), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT91), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n376_), .A2(new_n375_), .ZN(new_n390_));
  NOR4_X1   g189(.A1(new_n362_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT90), .B1(new_n371_), .B2(new_n372_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n366_), .A2(new_n368_), .B1(new_n363_), .B2(KEYINPUT3), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n389_), .B1(new_n395_), .B2(new_n386_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G127gat), .B(G134gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G113gat), .B(G120gat), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n388_), .A2(new_n396_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT100), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(KEYINPUT100), .A3(new_n400_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n406_), .A2(new_n377_), .A3(new_n387_), .A4(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n404_), .A3(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n403_), .A2(KEYINPUT4), .A3(new_n408_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n388_), .A2(new_n396_), .A3(new_n411_), .A4(new_n402_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n404_), .B(KEYINPUT101), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n361_), .B(new_n409_), .C1(new_n410_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT33), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n403_), .A2(KEYINPUT4), .A3(new_n408_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n413_), .A3(new_n412_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n361_), .A4(new_n409_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n403_), .A2(KEYINPUT104), .A3(new_n408_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT104), .B1(new_n403_), .B2(new_n408_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n413_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n412_), .A2(new_n404_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n361_), .B1(new_n417_), .B2(new_n424_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n416_), .A2(new_n420_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT19), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G169gat), .A2(G176gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G183gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT25), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT25), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G183gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT26), .B(G190gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n433_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT23), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT23), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(G183gat), .A3(G190gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT96), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT24), .ZN(new_n447_));
  INV_X1    g246(.A(G169gat), .ZN(new_n448_));
  INV_X1    g247(.A(G176gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n445_), .A2(new_n446_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n446_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n440_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT97), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n430_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G169gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n449_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n443_), .B1(G183gat), .B2(G190gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n444_), .A2(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n443_), .A2(KEYINPUT85), .A3(G183gat), .A4(G190gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G183gat), .A2(G190gat), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n455_), .B(new_n457_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n453_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G197gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT94), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT94), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G197gat), .ZN(new_n469_));
  INV_X1    g268(.A(G204gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT21), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(G197gat), .B2(G204gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G218gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(G211gat), .ZN(new_n476_));
  INV_X1    g275(.A(G211gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(G218gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G211gat), .B(G218gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(KEYINPUT95), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n474_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n467_), .A2(new_n469_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G204gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n466_), .A2(new_n470_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT21), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n479_), .A2(new_n480_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(KEYINPUT95), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n486_), .A2(KEYINPUT21), .A3(new_n487_), .ZN(new_n492_));
  OAI22_X1  g291(.A1(new_n484_), .A2(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT20), .B1(new_n465_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n434_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n445_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n431_), .B1(new_n456_), .B2(new_n449_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n450_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n460_), .A2(new_n461_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n442_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT26), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n438_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  AOI221_X4 g306(.A(KEYINPUT86), .B1(new_n499_), .B2(new_n500_), .C1(new_n503_), .C2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n502_), .A2(new_n442_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n501_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n507_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n500_), .A2(new_n499_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n509_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n493_), .B1(new_n508_), .B2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(KEYINPUT99), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT99), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n435_), .A2(new_n437_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n497_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT26), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n506_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n518_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n523_), .A2(new_n462_), .A3(new_n501_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n513_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT86), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n512_), .A2(new_n509_), .A3(new_n513_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n517_), .B1(new_n528_), .B2(new_n493_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n429_), .B(new_n495_), .C1(new_n516_), .C2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G8gat), .B(G36gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT18), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G64gat), .B(G92gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535_));
  INV_X1    g334(.A(new_n492_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n491_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n489_), .A2(new_n490_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT94), .B(G197gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n487_), .B1(new_n539_), .B2(new_n470_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n472_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n536_), .A2(new_n537_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n526_), .A2(new_n542_), .A3(new_n527_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT20), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n465_), .B2(new_n493_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n535_), .B1(new_n546_), .B2(new_n428_), .ZN(new_n547_));
  AOI211_X1 g346(.A(KEYINPUT98), .B(new_n429_), .C1(new_n543_), .C2(new_n545_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n530_), .B(new_n534_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n534_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n547_), .A2(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n515_), .A2(KEYINPUT99), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n528_), .A2(new_n517_), .A3(new_n493_), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n428_), .B(new_n494_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n550_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n426_), .A2(new_n549_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n534_), .A2(KEYINPUT32), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n530_), .B(new_n557_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n409_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n361_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n415_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n546_), .A2(new_n428_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n495_), .B1(new_n516_), .B2(new_n529_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n564_), .B2(new_n428_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n558_), .B(new_n562_), .C1(new_n557_), .C2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n556_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n388_), .A2(new_n396_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n569_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G78gat), .B(G106gat), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT29), .B1(new_n395_), .B2(new_n386_), .ZN(new_n577_));
  INV_X1    g376(.A(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(G228gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(G228gat), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT93), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n493_), .A2(new_n577_), .A3(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G22gat), .B(G50gat), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n388_), .A2(new_n396_), .A3(KEYINPUT29), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n588_), .A2(new_n493_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n585_), .B(new_n587_), .C1(new_n589_), .C2(new_n584_), .ZN(new_n590_));
  AOI211_X1 g389(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n388_), .C2(new_n396_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n574_), .B1(new_n571_), .B2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n584_), .B1(new_n588_), .B2(new_n493_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n585_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n586_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  AND4_X1   g394(.A1(new_n576_), .A2(new_n590_), .A3(new_n592_), .A4(new_n595_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n590_), .A2(new_n595_), .B1(new_n576_), .B2(new_n592_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n567_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT27), .ZN(new_n600_));
  INV_X1    g399(.A(new_n549_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n546_), .A2(new_n428_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT98), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n546_), .A2(new_n535_), .A3(new_n428_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n534_), .B1(new_n605_), .B2(new_n530_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n600_), .B1(new_n601_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n561_), .A2(new_n415_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n590_), .A2(new_n595_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n576_), .A2(new_n592_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n590_), .A2(new_n576_), .A3(new_n592_), .A4(new_n595_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n549_), .B(KEYINPUT27), .C1(new_n534_), .C2(new_n565_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n607_), .A2(new_n608_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n599_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G15gat), .B(G43gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G71gat), .B(G99gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(new_n402_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G227gat), .A2(G233gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT88), .Z(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n508_), .B2(new_n514_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT31), .ZN(new_n627_));
  INV_X1    g426(.A(new_n625_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n526_), .A2(new_n527_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n627_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n623_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n630_), .A3(new_n622_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n635_), .A2(new_n633_), .A3(new_n561_), .A4(new_n415_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n613_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n607_), .A2(new_n638_), .A3(new_n614_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT105), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n607_), .A2(new_n638_), .A3(new_n641_), .A4(new_n614_), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n616_), .A2(new_n636_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n297_), .A2(new_n303_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n304_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n249_), .A3(new_n305_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n647_), .B(new_n648_), .C1(new_n308_), .C2(new_n262_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n248_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n647_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n648_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT82), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT82), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n654_), .B(new_n648_), .C1(new_n650_), .C2(new_n647_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n649_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(G113gat), .B(G141gat), .Z(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT83), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G169gat), .B(G197gat), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n658_), .B(new_n659_), .Z(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n656_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n649_), .B(new_n660_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n265_), .A2(new_n344_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT12), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n265_), .A2(new_n344_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n269_), .A2(KEYINPUT12), .A3(new_n330_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n668_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n666_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(G120gat), .B(G148gat), .Z(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n676_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n668_), .A2(new_n667_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n245_), .A2(new_n350_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n330_), .A2(KEYINPUT12), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n684_), .B(new_n685_), .C1(new_n261_), .C2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n675_), .B(new_n681_), .C1(new_n687_), .C2(new_n673_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n683_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT13), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT13), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n683_), .A2(new_n691_), .A3(new_n688_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  NOR4_X1   g492(.A1(new_n354_), .A2(new_n643_), .A3(new_n665_), .A4(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n291_), .A3(new_n562_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n690_), .A2(new_n692_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n664_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(KEYINPUT106), .A3(new_n353_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702_));
  INV_X1    g501(.A(new_n353_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n699_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n283_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n643_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(new_n704_), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G1gat), .B1(new_n707_), .B2(new_n608_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n695_), .A2(new_n696_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n697_), .A2(new_n708_), .A3(new_n709_), .ZN(G1324gat));
  NAND2_X1  g509(.A1(new_n549_), .A2(KEYINPUT27), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n565_), .A2(new_n534_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT27), .B1(new_n555_), .B2(new_n549_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n694_), .A2(new_n292_), .A3(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT107), .ZN(new_n718_));
  OAI21_X1  g517(.A(G8gat), .B1(new_n707_), .B2(new_n715_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n720_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n718_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g523(.A(G15gat), .B1(new_n707_), .B2(new_n636_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n726_), .ZN(new_n728_));
  INV_X1    g527(.A(G15gat), .ZN(new_n729_));
  INV_X1    g528(.A(new_n636_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n694_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n727_), .A2(new_n728_), .A3(new_n731_), .ZN(G1326gat));
  OAI21_X1  g531(.A(G22gat), .B1(new_n707_), .B2(new_n598_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT42), .ZN(new_n734_));
  INV_X1    g533(.A(G22gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n694_), .A2(new_n735_), .A3(new_n613_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1327gat));
  NOR2_X1   g536(.A1(new_n643_), .A2(new_n665_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n353_), .A2(new_n283_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(new_n698_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G29gat), .B1(new_n741_), .B2(new_n562_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n643_), .A2(KEYINPUT43), .A3(new_n288_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n640_), .A2(new_n642_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n608_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n713_), .A2(new_n714_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n613_), .B1(new_n556_), .B2(new_n566_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n636_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n745_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n287_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n284_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n744_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n743_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n700_), .A2(new_n703_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n758_), .A2(new_n359_), .A3(new_n608_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n742_), .B1(new_n759_), .B2(new_n760_), .ZN(G1328gat));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n762_));
  INV_X1    g561(.A(G36gat), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n738_), .A2(new_n740_), .A3(new_n763_), .A4(new_n716_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT110), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n758_), .A2(new_n715_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n763_), .B1(new_n768_), .B2(new_n760_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n762_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n769_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n765_), .B(KEYINPUT45), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(KEYINPUT46), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(G1329gat));
  INV_X1    g573(.A(G43gat), .ZN(new_n775_));
  OR3_X1    g574(.A1(new_n758_), .A2(new_n775_), .A3(new_n636_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n760_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n741_), .A2(new_n730_), .ZN(new_n778_));
  OAI22_X1  g577(.A1(new_n776_), .A2(new_n777_), .B1(G43gat), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g579(.A(G50gat), .B1(new_n741_), .B2(new_n613_), .ZN(new_n781_));
  INV_X1    g580(.A(G50gat), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n758_), .A2(new_n782_), .A3(new_n598_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(new_n783_), .B2(new_n760_), .ZN(G1331gat));
  NAND2_X1  g583(.A1(new_n693_), .A2(new_n665_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(new_n354_), .A3(new_n643_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G57gat), .B1(new_n786_), .B2(new_n562_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n785_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(new_n706_), .A3(new_n353_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT111), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(G57gat), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n562_), .A2(KEYINPUT112), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(G57gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n787_), .B1(new_n790_), .B2(new_n794_), .ZN(G1332gat));
  INV_X1    g594(.A(G64gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n786_), .A2(new_n796_), .A3(new_n716_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT48), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n790_), .A2(new_n716_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G64gat), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT48), .B(new_n796_), .C1(new_n790_), .C2(new_n716_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(G1333gat));
  INV_X1    g601(.A(G71gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n786_), .A2(new_n803_), .A3(new_n730_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n790_), .A2(new_n730_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(G71gat), .ZN(new_n807_));
  AOI211_X1 g606(.A(KEYINPUT49), .B(new_n803_), .C1(new_n790_), .C2(new_n730_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(G1334gat));
  NAND3_X1  g608(.A1(new_n786_), .A2(new_n318_), .A3(new_n613_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n790_), .A2(new_n613_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(G78gat), .ZN(new_n813_));
  AOI211_X1 g612(.A(KEYINPUT50), .B(new_n318_), .C1(new_n790_), .C2(new_n613_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(G1335gat));
  NOR4_X1   g614(.A1(new_n785_), .A2(new_n643_), .A3(new_n353_), .A4(new_n283_), .ZN(new_n816_));
  INV_X1    g615(.A(G85gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n562_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT43), .B1(new_n643_), .B2(new_n288_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n750_), .A2(new_n744_), .A3(new_n753_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n785_), .A2(new_n353_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n562_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n818_), .B1(new_n824_), .B2(new_n817_), .ZN(G1336gat));
  AOI21_X1  g624(.A(G92gat), .B1(new_n816_), .B2(new_n716_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n716_), .A2(G92gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT113), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n823_), .B2(new_n828_), .ZN(G1337gat));
  NOR2_X1   g628(.A1(new_n636_), .A2(new_n218_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n816_), .A2(new_n830_), .B1(KEYINPUT114), .B2(KEYINPUT51), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n823_), .A2(new_n730_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n214_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n833_), .B(new_n834_), .Z(G1338gat));
  OAI211_X1 g634(.A(new_n613_), .B(new_n822_), .C1(new_n743_), .C2(new_n754_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n215_), .B1(new_n836_), .B2(KEYINPUT115), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n821_), .A2(new_n839_), .A3(new_n613_), .A4(new_n822_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n837_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n838_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n816_), .A2(new_n215_), .A3(new_n613_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n836_), .A2(KEYINPUT115), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(G106gat), .A3(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT116), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n848_), .B2(KEYINPUT52), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT53), .B1(new_n844_), .B2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n837_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(KEYINPUT52), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n842_), .A2(new_n843_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n845_), .A4(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n850_), .A2(new_n855_), .ZN(G1339gat));
  NAND4_X1  g655(.A1(new_n288_), .A2(new_n665_), .A3(new_n698_), .A4(new_n353_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n651_), .A2(new_n648_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n647_), .B(new_n652_), .C1(new_n308_), .C2(new_n262_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n661_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n663_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n864_), .A2(new_n688_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n671_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n672_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n669_), .A2(new_n670_), .A3(KEYINPUT55), .A4(new_n671_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT56), .B1(new_n870_), .B2(new_n682_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT56), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n872_), .B(new_n681_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n865_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n288_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n867_), .B1(new_n687_), .B2(new_n673_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n687_), .A2(new_n673_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n869_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n682_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n872_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n870_), .A2(KEYINPUT56), .A3(new_n682_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n884_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n865_), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT58), .B(new_n865_), .C1(new_n871_), .C2(new_n873_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n876_), .A2(new_n885_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n664_), .A2(new_n688_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n664_), .A2(new_n688_), .A3(KEYINPUT117), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n689_), .A2(new_n864_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n283_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  OAI221_X1 g699(.A(new_n283_), .B1(KEYINPUT118), .B2(KEYINPUT57), .C1(new_n895_), .C2(new_n897_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n889_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n859_), .B1(new_n902_), .B2(new_n703_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n716_), .A2(new_n608_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n730_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n903_), .A2(new_n613_), .A3(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G113gat), .B1(new_n906_), .B2(new_n664_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n902_), .A2(new_n703_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n859_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n905_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT59), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n912_), .A2(new_n598_), .A3(new_n913_), .A4(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n909_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n665_), .A2(KEYINPUT121), .ZN(new_n919_));
  MUX2_X1   g718(.A(KEYINPUT121), .B(new_n919_), .S(G113gat), .Z(new_n920_));
  AOI21_X1  g719(.A(new_n907_), .B1(new_n918_), .B2(new_n920_), .ZN(G1340gat));
  OAI211_X1 g720(.A(new_n916_), .B(new_n693_), .C1(new_n906_), .C2(new_n908_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(G120gat), .ZN(new_n923_));
  INV_X1    g722(.A(G120gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n698_), .B2(KEYINPUT60), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n906_), .B(new_n925_), .C1(KEYINPUT60), .C2(new_n924_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n923_), .A2(new_n926_), .ZN(G1341gat));
  AOI21_X1  g726(.A(G127gat), .B1(new_n906_), .B2(new_n353_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n353_), .A2(G127gat), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT122), .Z(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n918_), .B2(new_n930_), .ZN(G1342gat));
  OAI211_X1 g730(.A(new_n916_), .B(new_n753_), .C1(new_n906_), .C2(new_n908_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(G134gat), .ZN(new_n933_));
  INV_X1    g732(.A(G134gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n906_), .A2(new_n934_), .A3(new_n705_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1343gat));
  NOR4_X1   g735(.A1(new_n716_), .A2(new_n608_), .A3(new_n598_), .A4(new_n730_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n912_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n664_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g739(.A1(new_n912_), .A2(new_n937_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n698_), .ZN(new_n942_));
  XOR2_X1   g741(.A(KEYINPUT123), .B(G148gat), .Z(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1345gat));
  NOR2_X1   g743(.A1(new_n941_), .A2(new_n703_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT61), .B(G155gat), .Z(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1346gat));
  OR3_X1    g746(.A1(new_n941_), .A2(G162gat), .A3(new_n283_), .ZN(new_n948_));
  OAI21_X1  g747(.A(G162gat), .B1(new_n941_), .B2(new_n288_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1347gat));
  NOR2_X1   g749(.A1(new_n903_), .A2(new_n613_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n715_), .A2(new_n637_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  OAI211_X1 g752(.A(KEYINPUT62), .B(G169gat), .C1(new_n953_), .C2(new_n665_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n952_), .ZN(new_n955_));
  NOR4_X1   g754(.A1(new_n903_), .A2(new_n665_), .A3(new_n613_), .A4(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n456_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n958_), .B1(new_n956_), .B2(new_n448_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n954_), .A2(new_n957_), .A3(new_n959_), .ZN(G1348gat));
  OAI21_X1  g759(.A(new_n449_), .B1(new_n953_), .B2(new_n698_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n951_), .A2(KEYINPUT124), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n963_), .B1(new_n903_), .B2(new_n613_), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n698_), .A2(new_n955_), .A3(new_n449_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n962_), .A2(new_n964_), .A3(new_n965_), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n961_), .A2(new_n966_), .ZN(G1349gat));
  NOR3_X1   g766(.A1(new_n953_), .A2(new_n438_), .A3(new_n703_), .ZN(new_n968_));
  NAND4_X1  g767(.A1(new_n962_), .A2(new_n353_), .A3(new_n952_), .A4(new_n964_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n434_), .B2(new_n969_), .ZN(G1350gat));
  OAI21_X1  g769(.A(G190gat), .B1(new_n953_), .B2(new_n288_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n705_), .A2(new_n439_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n953_), .B2(new_n972_), .ZN(G1351gat));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n974_));
  NOR3_X1   g773(.A1(new_n715_), .A2(new_n746_), .A3(new_n730_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n912_), .A2(new_n974_), .A3(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(new_n975_), .ZN(new_n977_));
  OAI21_X1  g776(.A(KEYINPUT125), .B1(new_n903_), .B2(new_n977_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n976_), .A2(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(G197gat), .B1(new_n979_), .B2(new_n664_), .ZN(new_n980_));
  AOI211_X1 g779(.A(new_n466_), .B(new_n665_), .C1(new_n976_), .C2(new_n978_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n980_), .A2(new_n981_), .ZN(G1352gat));
  NOR2_X1   g781(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n983_));
  INV_X1    g782(.A(new_n983_), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n698_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n985_));
  AOI21_X1  g784(.A(new_n984_), .B1(new_n979_), .B2(new_n985_), .ZN(new_n986_));
  INV_X1    g785(.A(new_n985_), .ZN(new_n987_));
  AOI211_X1 g786(.A(new_n987_), .B(new_n983_), .C1(new_n976_), .C2(new_n978_), .ZN(new_n988_));
  NOR2_X1   g787(.A1(new_n986_), .A2(new_n988_), .ZN(G1353gat));
  NOR2_X1   g788(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n990_));
  INV_X1    g789(.A(new_n990_), .ZN(new_n991_));
  INV_X1    g790(.A(KEYINPUT63), .ZN(new_n992_));
  OAI21_X1  g791(.A(new_n353_), .B1(new_n992_), .B2(new_n477_), .ZN(new_n993_));
  XOR2_X1   g792(.A(new_n993_), .B(KEYINPUT127), .Z(new_n994_));
  INV_X1    g793(.A(new_n994_), .ZN(new_n995_));
  AOI21_X1  g794(.A(new_n991_), .B1(new_n979_), .B2(new_n995_), .ZN(new_n996_));
  AOI211_X1 g795(.A(new_n990_), .B(new_n994_), .C1(new_n976_), .C2(new_n978_), .ZN(new_n997_));
  NOR2_X1   g796(.A1(new_n996_), .A2(new_n997_), .ZN(G1354gat));
  NAND3_X1  g797(.A1(new_n979_), .A2(new_n475_), .A3(new_n705_), .ZN(new_n999_));
  AOI21_X1  g798(.A(new_n288_), .B1(new_n976_), .B2(new_n978_), .ZN(new_n1000_));
  OAI21_X1  g799(.A(new_n999_), .B1(new_n475_), .B2(new_n1000_), .ZN(G1355gat));
endmodule


