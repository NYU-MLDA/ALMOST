//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n955_, new_n956_, new_n957_, new_n959_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n982_, new_n983_,
    new_n984_, new_n986_, new_n987_, new_n989_, new_n990_, new_n992_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1002_, new_n1003_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT74), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OAI211_X1 g005(.A(KEYINPUT74), .B(KEYINPUT14), .C1(new_n202_), .C2(new_n203_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT75), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n211_), .A3(new_n207_), .A4(new_n208_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G1gat), .B(G8gat), .Z(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n210_), .A2(new_n214_), .A3(new_n212_), .ZN(new_n217_));
  INV_X1    g016(.A(G36gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G29gat), .ZN(new_n219_));
  INV_X1    g018(.A(G29gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G36gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT71), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G29gat), .B(G36gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT71), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G43gat), .B(G50gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n224_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n216_), .A2(new_n217_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n234_));
  OAI211_X1 g033(.A(G229gat), .B(G233gat), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n217_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n214_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n230_), .A2(KEYINPUT15), .A3(new_n231_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT15), .B1(new_n230_), .B2(new_n231_), .ZN(new_n239_));
  OAI22_X1  g038(.A1(new_n236_), .A2(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n216_), .A2(new_n217_), .A3(new_n232_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT77), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n235_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n235_), .B2(new_n244_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT24), .ZN(new_n252_));
  INV_X1    g051(.A(G169gat), .ZN(new_n253_));
  INV_X1    g052(.A(G176gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT79), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G190gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G183gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(new_n264_), .B2(G183gat), .ZN(new_n267_));
  INV_X1    g066(.A(G183gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n263_), .A2(new_n265_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n255_), .A2(new_n258_), .A3(KEYINPUT79), .A4(new_n259_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n253_), .A2(new_n254_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(KEYINPUT24), .A3(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n262_), .A2(new_n270_), .A3(new_n271_), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT22), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n254_), .B1(new_n276_), .B2(KEYINPUT80), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(new_n253_), .ZN(new_n278_));
  OR2_X1    g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n258_), .A2(new_n279_), .A3(new_n259_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285_));
  INV_X1    g084(.A(G15gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(G71gat), .ZN(new_n288_));
  INV_X1    g087(.A(G99gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n284_), .A2(new_n290_), .ZN(new_n293_));
  INV_X1    g092(.A(G134gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G127gat), .ZN(new_n295_));
  INV_X1    g094(.A(G127gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G134gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT82), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n301_));
  INV_X1    g100(.A(G120gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G113gat), .ZN(new_n303_));
  INV_X1    g102(.A(G113gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G120gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT83), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n308_));
  OAI22_X1  g107(.A1(new_n300_), .A2(new_n301_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n295_), .A2(new_n297_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT82), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n304_), .A2(G120gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n302_), .A2(G113gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT83), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n311_), .A2(new_n314_), .A3(new_n299_), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n309_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n292_), .A2(new_n293_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT81), .B(G43gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT31), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n318_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n293_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n317_), .B1(new_n326_), .B2(new_n291_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n325_), .B1(new_n327_), .B2(new_n319_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n268_), .A2(KEYINPUT25), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n265_), .A2(new_n334_), .A3(KEYINPUT92), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT92), .B1(new_n265_), .B2(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n263_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n274_), .A2(new_n258_), .A3(new_n259_), .A4(new_n255_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n253_), .A2(KEYINPUT22), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n276_), .A2(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT93), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n254_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n280_), .A2(new_n273_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n338_), .A2(new_n340_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G197gat), .ZN(new_n350_));
  INV_X1    g149(.A(G204gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT21), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G211gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n357_), .A2(G218gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT87), .B1(new_n357_), .B2(G218gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(KEYINPUT21), .A3(new_n353_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n356_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n352_), .A2(new_n353_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n363_), .B(KEYINPUT21), .C1(new_n358_), .C2(new_n359_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n333_), .B1(new_n349_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT94), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n364_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n282_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n282_), .B2(new_n368_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n332_), .B(new_n366_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n263_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n265_), .A2(new_n334_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n375_), .B2(new_n335_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n276_), .A2(G169gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n253_), .A2(KEYINPUT22), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT93), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n380_));
  AOI21_X1  g179(.A(G176gat), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OAI22_X1  g180(.A1(new_n376_), .A2(new_n339_), .B1(new_n381_), .B2(new_n347_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n368_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n365_), .A2(new_n281_), .A3(new_n275_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT20), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n331_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G8gat), .B(G36gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n371_), .A2(new_n386_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n333_), .B1(new_n382_), .B2(new_n368_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n393_), .A2(new_n332_), .A3(new_n384_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n366_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n331_), .B2(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT27), .B(new_n392_), .C1(new_n396_), .C2(new_n391_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n399_), .A2(G155gat), .A3(G162gat), .ZN(new_n400_));
  INV_X1    g199(.A(G155gat), .ZN(new_n401_));
  INV_X1    g200(.A(G162gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT85), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n398_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n408_));
  NAND3_X1  g207(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G141gat), .ZN(new_n411_));
  INV_X1    g210(.A(G148gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT3), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(G141gat), .B2(G148gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n405_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n413_), .A2(new_n415_), .B1(new_n416_), .B2(KEYINPUT2), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n404_), .B1(new_n410_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n411_), .A2(new_n412_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n407_), .A2(new_n409_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n398_), .A2(KEYINPUT1), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(G155gat), .A3(G162gat), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT85), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n399_), .B1(G155gat), .B2(G162gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n420_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n316_), .B(new_n309_), .C1(new_n418_), .C2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n413_), .A2(new_n415_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n416_), .A2(KEYINPUT2), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n410_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n425_), .A2(new_n426_), .B1(G155gat), .B2(G162gat), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n421_), .B(new_n423_), .C1(new_n400_), .C2(new_n403_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n420_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n432_), .A2(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n317_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n429_), .A2(new_n437_), .A3(KEYINPUT4), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n432_), .A2(new_n433_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n434_), .A2(new_n435_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n316_), .A4(new_n309_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n438_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n429_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G85gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT0), .B(G57gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(new_n452_), .A3(new_n447_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT27), .ZN(new_n457_));
  OAI211_X1 g256(.A(KEYINPUT20), .B(new_n332_), .C1(new_n382_), .C2(new_n368_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n282_), .A2(new_n368_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT94), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n282_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n332_), .B1(new_n393_), .B2(new_n384_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n391_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n391_), .B1(new_n371_), .B2(new_n386_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n457_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n397_), .A2(new_n456_), .A3(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G22gat), .B(G50gat), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT29), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n436_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n436_), .B2(new_n471_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n470_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n476_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n469_), .A3(new_n474_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n471_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n481_));
  OAI211_X1 g280(.A(G228gat), .B(G233gat), .C1(new_n481_), .C2(new_n365_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n483_), .B(new_n368_), .C1(new_n436_), .C2(new_n471_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G78gat), .B(G106gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT88), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n487_), .B1(new_n488_), .B2(KEYINPUT89), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n482_), .A2(new_n484_), .A3(new_n490_), .A4(new_n486_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n480_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT90), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n488_), .A2(KEYINPUT91), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n487_), .A2(new_n479_), .A3(new_n477_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n488_), .A2(KEYINPUT91), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n492_), .B2(KEYINPUT90), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n468_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n460_), .A2(new_n461_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n332_), .B1(new_n501_), .B2(new_n366_), .ZN(new_n502_));
  OAI211_X1 g301(.A(KEYINPUT32), .B(new_n391_), .C1(new_n502_), .C2(new_n394_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n454_), .A2(new_n455_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n458_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n501_), .A2(new_n505_), .B1(new_n331_), .B2(new_n385_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n391_), .A2(KEYINPUT32), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n506_), .A2(KEYINPUT99), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT99), .B1(new_n506_), .B2(new_n507_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n503_), .B(new_n504_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n455_), .A2(KEYINPUT33), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT33), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n446_), .A2(new_n512_), .A3(new_n452_), .A4(new_n447_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT98), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n429_), .A2(new_n437_), .A3(KEYINPUT4), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n445_), .A2(new_n439_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT97), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT97), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n438_), .A2(new_n519_), .A3(new_n439_), .A4(new_n445_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n429_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n453_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n515_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n525_));
  AOI211_X1 g324(.A(KEYINPUT98), .B(new_n523_), .C1(new_n518_), .C2(new_n520_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n514_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n528_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n464_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(KEYINPUT96), .A3(new_n392_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n510_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n489_), .A2(new_n491_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n477_), .A2(new_n479_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n493_), .A3(new_n498_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n329_), .B(new_n500_), .C1(new_n533_), .C2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n397_), .A2(new_n467_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n504_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n251_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G127gat), .B(G155gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT16), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G183gat), .B(G211gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G78gat), .ZN(new_n555_));
  INV_X1    g354(.A(G78gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n555_), .A2(new_n557_), .B1(KEYINPUT11), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(KEYINPUT11), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n555_), .A2(new_n557_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n216_), .A2(new_n217_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT76), .Z(new_n566_));
  OR2_X1    g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n566_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n563_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n551_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n549_), .B(KEYINPUT17), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n573_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G134gat), .B(G162gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  OR2_X1    g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT6), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n585_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT8), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT8), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n594_), .B(new_n585_), .C1(new_n588_), .C2(new_n591_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(G106gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT10), .B(G99gat), .Z(new_n598_));
  AOI21_X1  g397(.A(new_n591_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT65), .B(G92gat), .ZN(new_n600_));
  INV_X1    g399(.A(G85gat), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(KEYINPUT9), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT66), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n583_), .A2(KEYINPUT9), .A3(new_n584_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n604_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n599_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI22_X1  g408(.A1(new_n596_), .A2(new_n609_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n593_), .A2(new_n595_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n232_), .A3(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT34), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT35), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n612_), .B2(KEYINPUT72), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n613_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n617_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n610_), .A2(new_n612_), .A3(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n620_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n581_), .B(new_n582_), .C1(new_n622_), .C2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n612_), .A2(KEYINPUT72), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n618_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n628_), .A2(new_n612_), .A3(new_n610_), .A4(new_n623_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n629_), .A2(new_n580_), .A3(new_n579_), .A4(new_n621_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n626_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n576_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT5), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT70), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n603_), .A2(new_n605_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT66), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n645_), .A2(new_n599_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(KEYINPUT68), .A3(new_n562_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n611_), .A2(new_n562_), .A3(new_n608_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT68), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT69), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT69), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n647_), .A2(new_n650_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n611_), .A2(new_n608_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n563_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT64), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n648_), .A2(new_n659_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n646_), .A2(KEYINPUT12), .A3(new_n562_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT12), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n655_), .B2(new_n563_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n641_), .B1(new_n661_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n666_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n655_), .A2(new_n665_), .A3(new_n563_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n662_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n640_), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n671_), .B(new_n672_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT13), .B1(new_n668_), .B2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n661_), .A2(new_n667_), .A3(new_n640_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT13), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n671_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n675_), .B(new_n676_), .C1(new_n677_), .C2(new_n641_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n636_), .B1(new_n674_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n545_), .A2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT100), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n202_), .A3(new_n504_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT38), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n684_), .A2(KEYINPUT101), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(KEYINPUT101), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n674_), .A2(new_n678_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n572_), .A2(new_n575_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n688_), .A2(new_n251_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n626_), .A2(new_n630_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n202_), .B1(new_n695_), .B2(new_n504_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n682_), .B1(new_n683_), .B2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n685_), .A2(new_n686_), .A3(new_n697_), .ZN(G1324gat));
  OAI21_X1  g497(.A(G8gat), .B1(new_n694_), .B2(new_n542_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT39), .ZN(new_n700_));
  INV_X1    g499(.A(new_n542_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n681_), .A2(new_n203_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g503(.A(G15gat), .B1(new_n694_), .B2(new_n329_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n708_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n329_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n681_), .A2(new_n286_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n713_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n709_), .A2(new_n710_), .A3(new_n714_), .A4(new_n715_), .ZN(G1326gat));
  OAI21_X1  g515(.A(G22gat), .B1(new_n694_), .B2(new_n541_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT105), .Z(new_n718_));
  OR2_X1    g517(.A1(new_n718_), .A2(KEYINPUT42), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(KEYINPUT42), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n541_), .A2(G22gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT106), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n681_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n719_), .A2(new_n720_), .A3(new_n723_), .ZN(G1327gat));
  NOR2_X1   g523(.A1(new_n576_), .A2(new_n691_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n687_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n545_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G29gat), .B1(new_n728_), .B2(new_n504_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n540_), .A2(new_n544_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n633_), .A2(new_n635_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(KEYINPUT43), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735_));
  INV_X1    g534(.A(new_n635_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n626_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT107), .B1(new_n633_), .B2(new_n635_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n730_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n735_), .B1(new_n742_), .B2(KEYINPUT43), .ZN(new_n743_));
  AOI22_X1  g542(.A1(new_n540_), .A2(new_n544_), .B1(new_n740_), .B2(new_n739_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n744_), .A2(KEYINPUT108), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n734_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n251_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n687_), .A2(new_n748_), .A3(new_n689_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(KEYINPUT44), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n742_), .A2(new_n735_), .A3(KEYINPUT43), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT108), .B1(new_n744_), .B2(new_n745_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n749_), .B1(new_n756_), .B2(new_n734_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n753_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n747_), .A2(new_n750_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n759_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n456_), .A2(new_n220_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n729_), .B1(new_n763_), .B2(new_n764_), .ZN(G1328gat));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n701_), .B1(new_n757_), .B2(KEYINPUT44), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n218_), .B1(new_n759_), .B2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n728_), .A2(new_n218_), .A3(new_n701_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT45), .Z(new_n771_));
  OAI21_X1  g570(.A(new_n766_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n771_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n767_), .B1(new_n753_), .B2(new_n758_), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT46), .B(new_n773_), .C1(new_n774_), .C2(new_n218_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n775_), .ZN(G1329gat));
  INV_X1    g575(.A(G43gat), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n329_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT109), .B1(new_n757_), .B2(KEYINPUT44), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n754_), .A2(new_n755_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n780_));
  NOR4_X1   g579(.A1(new_n780_), .A2(new_n752_), .A3(new_n761_), .A4(new_n749_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n762_), .B(new_n778_), .C1(new_n779_), .C2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(new_n727_), .B2(new_n329_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1330gat));
  OR3_X1    g586(.A1(new_n727_), .A2(G50gat), .A3(new_n541_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n541_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n790_), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT111), .B1(new_n790_), .B2(G50gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(G1331gat));
  NOR2_X1   g592(.A1(new_n687_), .A2(new_n748_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n693_), .A2(new_n576_), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(G57gat), .B1(new_n795_), .B2(new_n456_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n794_), .A2(new_n730_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n689_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n456_), .A2(G57gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(G1332gat));
  OAI21_X1  g600(.A(G64gat), .B1(new_n795_), .B2(new_n542_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT48), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n542_), .A2(G64gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n799_), .B2(new_n804_), .ZN(G1333gat));
  OAI21_X1  g604(.A(G71gat), .B1(new_n795_), .B2(new_n329_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT49), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n329_), .A2(G71gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n799_), .B2(new_n808_), .ZN(G1334gat));
  OAI21_X1  g608(.A(G78gat), .B1(new_n795_), .B2(new_n541_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT50), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n539_), .A2(new_n556_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n799_), .B2(new_n812_), .ZN(G1335gat));
  NAND2_X1  g612(.A1(new_n797_), .A2(new_n725_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT112), .ZN(new_n815_));
  AOI21_X1  g614(.A(G85gat), .B1(new_n815_), .B2(new_n504_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT113), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n794_), .A2(new_n689_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n780_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n456_), .A2(new_n601_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n817_), .B1(new_n819_), .B2(new_n820_), .ZN(G1336gat));
  AOI21_X1  g620(.A(G92gat), .B1(new_n815_), .B2(new_n701_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n701_), .A2(new_n600_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n819_), .B2(new_n823_), .ZN(G1337gat));
  AND2_X1   g623(.A1(new_n711_), .A2(new_n598_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n815_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT114), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n289_), .B1(new_n819_), .B2(new_n711_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1338gat));
  NAND3_X1  g630(.A1(new_n815_), .A2(new_n597_), .A3(new_n539_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n819_), .A2(new_n539_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(G106gat), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT52), .B(new_n597_), .C1(new_n819_), .C2(new_n539_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT53), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n832_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1339gat));
  NOR2_X1   g640(.A1(new_n251_), .A2(new_n304_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n664_), .A2(new_n666_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n660_), .B1(new_n845_), .B2(new_n651_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n667_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n663_), .B(KEYINPUT55), .C1(new_n664_), .C2(new_n666_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n641_), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n844_), .B(KEYINPUT56), .C1(new_n850_), .C2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n243_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n243_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n240_), .A2(new_n241_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n247_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n248_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT116), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n248_), .A2(new_n860_), .A3(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n675_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n852_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n850_), .B2(new_n851_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n850_), .A2(KEYINPUT56), .A3(new_n851_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n844_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT58), .B1(new_n864_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n843_), .B1(new_n869_), .B2(new_n732_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n864_), .A2(new_n868_), .A3(KEYINPUT58), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872_));
  INV_X1    g671(.A(new_n867_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n873_), .A2(new_n865_), .A3(KEYINPUT118), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n865_), .A2(KEYINPUT118), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n677_), .A2(new_n640_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n872_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(KEYINPUT119), .A3(new_n731_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n870_), .A2(new_n871_), .A3(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n862_), .B1(new_n668_), .B2(new_n673_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT117), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n748_), .B(new_n675_), .C1(new_n873_), .C2(new_n865_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n884_), .B(new_n862_), .C1(new_n668_), .C2(new_n673_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(new_n883_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n692_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n887_), .A2(new_n888_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n886_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n689_), .B1(new_n880_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n679_), .B2(new_n251_), .ZN(new_n899_));
  AND4_X1   g698(.A1(new_n898_), .A2(new_n687_), .A3(new_n251_), .A4(new_n798_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n679_), .A2(new_n898_), .A3(new_n251_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n687_), .A2(new_n798_), .A3(new_n251_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT115), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n904_), .A3(KEYINPUT54), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n901_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n896_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n701_), .A2(new_n539_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n711_), .A3(new_n504_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(KEYINPUT59), .B1(new_n908_), .B2(new_n911_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n886_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n891_), .B1(new_n886_), .B2(new_n889_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n870_), .A2(new_n871_), .A3(new_n879_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n576_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(KEYINPUT59), .B(new_n911_), .C1(new_n917_), .C2(new_n906_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n842_), .B1(new_n912_), .B2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n908_), .A2(new_n911_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n304_), .B1(new_n922_), .B2(new_n251_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(new_n921_), .A3(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n842_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n915_), .A2(new_n916_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n906_), .B1(new_n927_), .B2(new_n689_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n928_), .B2(new_n910_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n925_), .B1(new_n929_), .B2(new_n918_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n910_), .ZN(new_n931_));
  AOI21_X1  g730(.A(G113gat), .B1(new_n931_), .B2(new_n748_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT121), .B1(new_n930_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n924_), .A2(new_n933_), .ZN(G1340gat));
  AOI21_X1  g733(.A(new_n687_), .B1(new_n929_), .B2(new_n918_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT122), .B(G120gat), .Z(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n687_), .B2(KEYINPUT60), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(KEYINPUT60), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(KEYINPUT123), .B2(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n939_), .B1(KEYINPUT123), .B2(new_n937_), .ZN(new_n940_));
  OAI22_X1  g739(.A1(new_n935_), .A2(new_n936_), .B1(new_n922_), .B2(new_n940_), .ZN(G1341gat));
  NOR2_X1   g740(.A1(new_n689_), .A2(new_n296_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n912_), .B2(new_n919_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n296_), .B1(new_n922_), .B2(new_n689_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n942_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(new_n929_), .B2(new_n918_), .ZN(new_n948_));
  AOI21_X1  g747(.A(G127gat), .B1(new_n931_), .B2(new_n576_), .ZN(new_n949_));
  OAI21_X1  g748(.A(KEYINPUT124), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n946_), .A2(new_n950_), .ZN(G1342gat));
  NAND3_X1  g750(.A1(new_n931_), .A2(new_n294_), .A3(new_n692_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n732_), .B1(new_n929_), .B2(new_n918_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(new_n294_), .ZN(G1343gat));
  NOR3_X1   g753(.A1(new_n711_), .A2(new_n701_), .A3(new_n456_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n908_), .A2(new_n539_), .A3(new_n955_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n956_), .A2(new_n251_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(new_n411_), .ZN(G1344gat));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n687_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(new_n412_), .ZN(G1345gat));
  NOR2_X1   g759(.A1(new_n956_), .A2(new_n689_), .ZN(new_n961_));
  XOR2_X1   g760(.A(KEYINPUT61), .B(G155gat), .Z(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n962_), .ZN(G1346gat));
  INV_X1    g762(.A(new_n956_), .ZN(new_n964_));
  AOI21_X1  g763(.A(G162gat), .B1(new_n964_), .B2(new_n692_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n402_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n964_), .B2(new_n966_), .ZN(G1347gat));
  AOI21_X1  g766(.A(new_n253_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n542_), .A2(new_n504_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n969_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n970_), .A2(new_n539_), .A3(new_n329_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n908_), .A2(new_n971_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n968_), .B1(new_n972_), .B2(new_n251_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n972_), .ZN(new_n976_));
  OAI211_X1 g775(.A(new_n976_), .B(new_n748_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n977_));
  OAI221_X1 g776(.A(new_n968_), .B1(KEYINPUT125), .B2(KEYINPUT62), .C1(new_n972_), .C2(new_n251_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n975_), .A2(new_n977_), .A3(new_n978_), .ZN(G1348gat));
  NAND2_X1  g778(.A1(new_n976_), .A2(new_n688_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(new_n980_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g780(.A1(new_n976_), .A2(new_n576_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(G183gat), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n336_), .A2(new_n337_), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n983_), .B1(new_n984_), .B2(new_n982_), .ZN(G1350gat));
  OAI21_X1  g784(.A(G190gat), .B1(new_n972_), .B2(new_n732_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n692_), .A2(new_n263_), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n986_), .B1(new_n972_), .B2(new_n987_), .ZN(G1351gat));
  NAND4_X1  g787(.A1(new_n908_), .A2(new_n539_), .A3(new_n329_), .A4(new_n969_), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n989_), .A2(new_n251_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n990_), .B(new_n350_), .ZN(G1352gat));
  NOR2_X1   g790(.A1(new_n989_), .A2(new_n687_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(new_n351_), .ZN(G1353gat));
  AOI21_X1  g792(.A(new_n689_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n994_));
  INV_X1    g793(.A(new_n994_), .ZN(new_n995_));
  NOR2_X1   g794(.A1(new_n989_), .A2(new_n995_), .ZN(new_n996_));
  NOR2_X1   g795(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n997_));
  XNOR2_X1  g796(.A(new_n997_), .B(KEYINPUT126), .ZN(new_n998_));
  XNOR2_X1  g797(.A(new_n998_), .B(KEYINPUT127), .ZN(new_n999_));
  INV_X1    g798(.A(new_n999_), .ZN(new_n1000_));
  XNOR2_X1  g799(.A(new_n996_), .B(new_n1000_), .ZN(G1354gat));
  OAI21_X1  g800(.A(G218gat), .B1(new_n989_), .B2(new_n732_), .ZN(new_n1002_));
  OR2_X1    g801(.A1(new_n691_), .A2(G218gat), .ZN(new_n1003_));
  OAI21_X1  g802(.A(new_n1002_), .B1(new_n989_), .B2(new_n1003_), .ZN(G1355gat));
endmodule


