//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202_));
  OR2_X1    g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT90), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT90), .B1(new_n206_), .B2(new_n207_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT2), .ZN(new_n214_));
  OR2_X1    g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n213_), .A2(new_n214_), .B1(KEYINPUT3), .B2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n205_), .B1(new_n211_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n204_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n206_), .B(KEYINPUT89), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n203_), .A2(new_n218_), .A3(new_n204_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n202_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(new_n214_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n210_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n215_), .A2(KEYINPUT3), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .A4(new_n208_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n205_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(KEYINPUT91), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n224_), .A2(new_n232_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(KEYINPUT100), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n217_), .A2(new_n223_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT100), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n239_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G57gat), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT103), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G1gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT102), .B(KEYINPUT0), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G29gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n249_), .B(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n239_), .A2(KEYINPUT4), .A3(new_n244_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n224_), .A2(new_n232_), .A3(new_n254_), .A4(new_n238_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n245_), .B(KEYINPUT101), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n246_), .B(new_n252_), .C1(new_n253_), .C2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT33), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n239_), .A2(new_n244_), .A3(KEYINPUT4), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT33), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n246_), .A4(new_n252_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n239_), .A2(new_n244_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n264_), .A2(KEYINPUT104), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(KEYINPUT104), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n256_), .A3(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n255_), .A2(new_n245_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n252_), .B1(new_n268_), .B2(new_n260_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n259_), .A2(new_n263_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G8gat), .B(G36gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT18), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT98), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT20), .ZN(new_n277_));
  INV_X1    g076(.A(G169gat), .ZN(new_n278_));
  INV_X1    g077(.A(G176gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(KEYINPUT24), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT25), .B(G183gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G190gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G183gat), .ZN(new_n286_));
  INV_X1    g085(.A(G190gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT23), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(G183gat), .A3(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT96), .ZN(new_n292_));
  OR3_X1    g091(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n282_), .B(new_n285_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n281_), .B(KEYINPUT97), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT22), .B(G169gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n279_), .B2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n289_), .B1(G183gat), .B2(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n290_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n289_), .A2(KEYINPUT85), .A3(G183gat), .A4(G190gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n299_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n296_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G211gat), .B(G218gat), .Z(new_n308_));
  INV_X1    g107(.A(KEYINPUT95), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT95), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT94), .B(G197gat), .ZN(new_n313_));
  INV_X1    g112(.A(G204gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(G197gat), .B2(G204gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n310_), .A2(new_n312_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G197gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n314_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n316_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n321_), .A2(new_n316_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n311_), .B(new_n309_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n277_), .B1(new_n307_), .B2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(KEYINPUT25), .B(G183gat), .Z(new_n329_));
  NAND2_X1  g128(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT26), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n329_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n282_), .A2(new_n293_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n336_), .A2(new_n304_), .A3(new_n337_), .ZN(new_n338_));
  OR3_X1    g137(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT84), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n287_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n286_), .A3(new_n330_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n291_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT86), .B1(new_n338_), .B2(new_n345_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n318_), .A2(new_n322_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n304_), .A2(new_n337_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n343_), .B2(new_n330_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n283_), .B1(new_n350_), .B2(new_n334_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT86), .ZN(new_n353_));
  INV_X1    g152(.A(new_n345_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n346_), .A2(new_n347_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n328_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n276_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  AOI211_X1 g160(.A(KEYINPUT98), .B(new_n361_), .C1(new_n328_), .C2(new_n356_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT20), .B1(new_n307_), .B2(new_n327_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n346_), .A2(new_n355_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(new_n327_), .ZN(new_n368_));
  AOI211_X1 g167(.A(KEYINPUT99), .B(new_n347_), .C1(new_n346_), .C2(new_n355_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n361_), .B(new_n365_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n275_), .B1(new_n363_), .B2(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n370_), .B(new_n274_), .C1(new_n360_), .C2(new_n362_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n270_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n261_), .A2(new_n246_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n252_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n258_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n274_), .A2(KEYINPUT32), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n370_), .B(new_n379_), .C1(new_n360_), .C2(new_n362_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n357_), .A2(new_n359_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n365_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n359_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n378_), .B(new_n380_), .C1(new_n383_), .C2(new_n379_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n374_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(G228gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(G228gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT93), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n327_), .B(new_n392_), .C1(new_n241_), .C2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G22gat), .B(G50gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n224_), .A2(new_n232_), .A3(KEYINPUT29), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n397_), .A2(new_n327_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n394_), .B(new_n396_), .C1(new_n398_), .C2(new_n392_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n392_), .B1(new_n397_), .B2(new_n327_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n394_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n395_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n224_), .A2(new_n232_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n405_), .B2(new_n393_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n404_), .A3(new_n393_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  AOI211_X1 g210(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n224_), .C2(new_n232_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n409_), .B1(new_n406_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n403_), .A2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n399_), .A2(new_n411_), .A3(new_n402_), .A4(new_n413_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n385_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT27), .ZN(new_n420_));
  INV_X1    g219(.A(new_n360_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n357_), .A2(new_n276_), .A3(new_n359_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n274_), .B1(new_n423_), .B2(new_n370_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n373_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n420_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n378_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n373_), .B(KEYINPUT27), .C1(new_n383_), .C2(new_n274_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n417_), .A4(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n419_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT31), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT88), .Z(new_n433_));
  NOR3_X1   g232(.A1(new_n338_), .A2(KEYINPUT86), .A3(new_n345_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n353_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n433_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n346_), .A2(new_n355_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n431_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n438_), .A3(new_n431_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G15gat), .B(G43gat), .Z(new_n442_));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(KEYINPUT87), .B(KEYINPUT30), .Z(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(new_n238_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n436_), .A2(new_n438_), .A3(new_n431_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n439_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n377_), .A2(new_n448_), .A3(new_n258_), .A4(new_n451_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n417_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n426_), .A2(new_n428_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT105), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT105), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n426_), .A2(new_n454_), .A3(new_n457_), .A4(new_n428_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n430_), .A2(new_n452_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT9), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT64), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n464_));
  OAI22_X1  g263(.A1(new_n462_), .A2(KEYINPUT65), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n466_));
  INV_X1    g265(.A(G85gat), .ZN(new_n467_));
  INV_X1    g266(.A(G92gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT65), .B1(new_n470_), .B2(new_n462_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT10), .B(G99gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(G106gat), .B2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G99gat), .ZN(new_n481_));
  INV_X1    g280(.A(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n474_), .A2(new_n475_), .B1(KEYINPUT7), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n484_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT69), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT69), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n495_), .B(new_n484_), .C1(new_n491_), .C2(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n469_), .A2(new_n460_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT70), .B(KEYINPUT8), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n483_), .A2(KEYINPUT7), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n476_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n487_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n490_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT68), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n502_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT8), .B1(new_n508_), .B2(new_n497_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n500_), .A2(KEYINPUT73), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT73), .B1(new_n500_), .B2(new_n509_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n480_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT71), .B(G71gat), .Z(new_n513_));
  INV_X1    g312(.A(G78gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT71), .B(G71gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(G78gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n517_), .B(new_n515_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT12), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n512_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(KEYINPUT72), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT72), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n499_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n493_), .B2(KEYINPUT69), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n493_), .A2(new_n460_), .A3(new_n469_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n533_), .A2(new_n496_), .B1(new_n534_), .B2(KEYINPUT8), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n529_), .B(new_n531_), .C1(new_n535_), .C2(new_n479_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n499_), .B1(new_n508_), .B2(new_n495_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n496_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n509_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n529_), .A2(new_n531_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n539_), .A2(new_n480_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n536_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n528_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n479_), .B1(new_n500_), .B2(new_n509_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(new_n540_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n548_), .B2(new_n541_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G120gat), .B(G148gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G176gat), .B(G204gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n545_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT13), .ZN(new_n559_));
  OR3_X1    g358(.A1(new_n556_), .A2(KEYINPUT13), .A3(new_n557_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G29gat), .B(G36gat), .Z(new_n562_));
  XOR2_X1   g361(.A(G43gat), .B(G50gat), .Z(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT15), .Z(new_n565_));
  AND2_X1   g364(.A1(G15gat), .A2(G22gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(G15gat), .A2(G22gat), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G1gat), .A2(G8gat), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n569_), .A2(KEYINPUT14), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n568_), .A2(new_n570_), .A3(KEYINPUT78), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT78), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(KEYINPUT14), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT79), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT78), .B1(new_n568_), .B2(new_n570_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n573_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G1gat), .B(G8gat), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n576_), .A2(new_n582_), .A3(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n565_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n564_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n584_), .A2(new_n588_), .A3(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n576_), .A2(new_n582_), .A3(new_n580_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n582_), .B1(new_n576_), .B2(new_n580_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n564_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n589_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n590_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT82), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT82), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n598_), .B(new_n590_), .C1(new_n594_), .C2(new_n589_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n591_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G113gat), .B(G141gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT83), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n591_), .B(new_n604_), .C1(new_n597_), .C2(new_n599_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n459_), .A2(new_n561_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n547_), .A2(new_n588_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT73), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n539_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n500_), .A2(KEYINPUT73), .A3(new_n509_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n479_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n565_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n611_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n618_));
  NAND2_X1  g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n620_), .B(KEYINPUT35), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n611_), .B(new_n628_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n623_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT76), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT76), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n623_), .A2(new_n632_), .A3(new_n627_), .A4(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n623_), .A2(new_n629_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n626_), .B(KEYINPUT36), .Z(new_n635_));
  AOI22_X1  g434(.A1(new_n631_), .A2(new_n633_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n636_), .B(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(G231gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n586_), .B1(new_n640_), .B2(new_n386_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n584_), .A2(G231gat), .A3(G233gat), .A4(new_n585_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(new_n525_), .ZN(new_n644_));
  XOR2_X1   g443(.A(G127gat), .B(G155gat), .Z(new_n645_));
  XNOR2_X1  g444(.A(G183gat), .B(G211gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT17), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n644_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT81), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n644_), .A2(new_n530_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n644_), .A2(new_n530_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n649_), .A2(KEYINPUT17), .ZN(new_n655_));
  NOR4_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n650_), .A4(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n639_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n610_), .A2(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n660_), .A2(G1gat), .A3(new_n427_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT38), .Z(new_n662_));
  NOR3_X1   g461(.A1(new_n561_), .A2(new_n658_), .A3(new_n609_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT106), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT106), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n459_), .A2(new_n636_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G1gat), .B1(new_n667_), .B2(new_n427_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n662_), .A2(new_n668_), .ZN(G1324gat));
  INV_X1    g468(.A(new_n428_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT27), .B1(new_n372_), .B2(new_n373_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G8gat), .B1(new_n667_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n660_), .A2(G8gat), .A3(new_n672_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(new_n674_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n675_), .A2(new_n678_), .A3(KEYINPUT40), .A4(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1325gat));
  OAI21_X1  g483(.A(G15gat), .B1(new_n667_), .B2(new_n452_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n660_), .A2(G15gat), .A3(new_n452_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(G1326gat));
  OAI21_X1  g489(.A(G22gat), .B1(new_n667_), .B2(new_n418_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT42), .Z(new_n692_));
  NOR3_X1   g491(.A1(new_n660_), .A2(G22gat), .A3(new_n418_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n631_), .A2(new_n633_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n634_), .A2(new_n635_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n657_), .A2(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n610_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G29gat), .B1(new_n699_), .B2(new_n378_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n638_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n636_), .A2(new_n637_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n459_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n456_), .A2(new_n458_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n417_), .A2(new_n427_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n670_), .A2(new_n671_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n417_), .B1(new_n374_), .B2(new_n384_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n452_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n639_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n704_), .A2(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n561_), .A2(new_n609_), .A3(new_n657_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(KEYINPUT44), .A3(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT44), .B1(new_n713_), .B2(new_n714_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n378_), .A2(G29gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n700_), .B1(new_n717_), .B2(new_n718_), .ZN(G1328gat));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n672_), .A2(G36gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n699_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n610_), .A2(new_n698_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n721_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT110), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT45), .ZN(new_n727_));
  INV_X1    g526(.A(G36gat), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n715_), .A2(new_n716_), .A3(new_n672_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n727_), .B(KEYINPUT46), .C1(new_n728_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n726_), .B(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n729_), .A2(new_n728_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n730_), .A2(new_n735_), .ZN(G1329gat));
  INV_X1    g535(.A(new_n452_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G43gat), .B1(new_n699_), .B2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n737_), .A2(G43gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n717_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n699_), .B2(new_n417_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n417_), .A2(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n717_), .B2(new_n743_), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n561_), .A2(new_n609_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(new_n459_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(new_n659_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G57gat), .B1(new_n747_), .B2(new_n378_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n666_), .A2(new_n609_), .A3(new_n561_), .A4(new_n657_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT111), .ZN(new_n750_));
  INV_X1    g549(.A(G57gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n378_), .B2(KEYINPUT112), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(KEYINPUT112), .B2(new_n751_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n748_), .B1(new_n750_), .B2(new_n753_), .ZN(G1332gat));
  INV_X1    g553(.A(G64gat), .ZN(new_n755_));
  INV_X1    g554(.A(new_n672_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n747_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n756_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G64gat), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT48), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT48), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n747_), .A2(new_n763_), .A3(new_n737_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n750_), .A2(new_n737_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G71gat), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT49), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT49), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1334gat));
  NAND3_X1  g568(.A1(new_n747_), .A2(new_n514_), .A3(new_n417_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n750_), .A2(new_n417_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G78gat), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT50), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(KEYINPUT50), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1335gat));
  NAND3_X1  g574(.A1(new_n561_), .A2(new_n609_), .A3(new_n658_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n704_), .B2(new_n712_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778_), .B2(new_n427_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n746_), .A2(new_n698_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n467_), .A3(new_n378_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1336gat));
  AOI21_X1  g581(.A(G92gat), .B1(new_n780_), .B2(new_n756_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n756_), .A2(G92gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT113), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n777_), .B2(new_n785_), .ZN(G1337gat));
  OAI21_X1  g585(.A(G99gat), .B1(new_n778_), .B2(new_n452_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n452_), .A2(new_n477_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n780_), .A2(new_n788_), .B1(KEYINPUT114), .B2(KEYINPUT51), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n790_), .B(new_n791_), .Z(G1338gat));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  INV_X1    g592(.A(new_n776_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n713_), .A2(new_n793_), .A3(new_n417_), .A4(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G106gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n793_), .B1(new_n777_), .B2(new_n417_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT116), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n713_), .A2(new_n417_), .A3(new_n794_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT115), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(G106gat), .A4(new_n795_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n798_), .A2(KEYINPUT52), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT116), .B(new_n804_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n780_), .A2(new_n482_), .A3(new_n417_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT53), .B1(new_n803_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n798_), .A2(KEYINPUT52), .A3(new_n802_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n805_), .A4(new_n806_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n604_), .B1(new_n595_), .B2(new_n590_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n587_), .A2(new_n589_), .A3(new_n596_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n607_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n556_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n544_), .B1(new_n528_), .B2(new_n543_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n545_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n528_), .A2(new_n543_), .A3(KEYINPUT55), .A4(new_n544_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n554_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n826_), .B(new_n554_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n818_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n813_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n542_), .B1(new_n547_), .B2(new_n540_), .ZN(new_n831_));
  OAI22_X1  g630(.A1(new_n615_), .A2(new_n526_), .B1(new_n831_), .B2(new_n548_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n820_), .B1(new_n832_), .B2(new_n546_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n545_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n822_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n824_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n826_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n824_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n840_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n818_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n828_), .A2(new_n829_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n830_), .A2(new_n841_), .A3(new_n639_), .A4(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n608_), .A2(new_n555_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n608_), .A2(new_n555_), .A3(KEYINPUT117), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n817_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n558_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n697_), .B1(new_n849_), .B2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n608_), .A2(new_n555_), .A3(KEYINPUT117), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT117), .B1(new_n608_), .B2(new_n555_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n851_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n854_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n697_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n843_), .A2(new_n855_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n658_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n559_), .A2(new_n560_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n703_), .A2(new_n609_), .A3(new_n865_), .A4(new_n657_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT54), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n756_), .A2(new_n427_), .A3(new_n452_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n418_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871_), .B2(new_n608_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n417_), .B1(new_n864_), .B2(new_n867_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(KEYINPUT120), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n869_), .A3(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n874_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n609_), .A2(KEYINPUT121), .ZN(new_n881_));
  MUX2_X1   g680(.A(KEYINPUT121), .B(new_n881_), .S(G113gat), .Z(new_n882_));
  AOI21_X1  g681(.A(new_n872_), .B1(new_n880_), .B2(new_n882_), .ZN(G1340gat));
  NAND3_X1  g682(.A1(new_n874_), .A2(new_n561_), .A3(new_n879_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G120gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n865_), .A2(KEYINPUT60), .ZN(new_n886_));
  MUX2_X1   g685(.A(new_n886_), .B(KEYINPUT60), .S(G120gat), .Z(new_n887_));
  NAND2_X1  g686(.A1(new_n871_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n888_), .ZN(G1341gat));
  AOI21_X1  g688(.A(G127gat), .B1(new_n871_), .B2(new_n657_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n657_), .A2(G127gat), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n891_), .B(KEYINPUT122), .Z(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n880_), .B2(new_n892_), .ZN(G1342gat));
  NAND3_X1  g692(.A1(new_n874_), .A2(new_n639_), .A3(new_n879_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G134gat), .ZN(new_n895_));
  OR3_X1    g694(.A1(new_n870_), .A2(G134gat), .A3(new_n697_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1343gat));
  NAND4_X1  g696(.A1(new_n672_), .A2(new_n378_), .A3(new_n417_), .A4(new_n452_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n864_), .B2(new_n867_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n608_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n561_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT123), .B(G148gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1345gat));
  NAND2_X1  g703(.A1(new_n899_), .A2(new_n657_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT61), .B(G155gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1346gat));
  INV_X1    g706(.A(G162gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n899_), .A2(new_n908_), .A3(new_n636_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n899_), .A2(new_n639_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n908_), .ZN(G1347gat));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n868_), .A2(new_n756_), .A3(new_n454_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n609_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n914_), .B2(new_n278_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n298_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT62), .B(G169gat), .C1(new_n913_), .C2(new_n609_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(G1348gat));
  INV_X1    g717(.A(new_n913_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G176gat), .B1(new_n919_), .B2(new_n561_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n865_), .A2(new_n279_), .A3(new_n672_), .A4(new_n453_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n920_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NOR3_X1   g724(.A1(new_n913_), .A2(new_n658_), .A3(new_n283_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n672_), .A2(new_n453_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n921_), .A2(new_n657_), .A3(new_n922_), .A4(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n928_), .B2(new_n286_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n913_), .B2(new_n703_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n636_), .A2(new_n284_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n913_), .B2(new_n931_), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n706_), .A2(new_n737_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n861_), .B1(new_n860_), .B2(new_n697_), .ZN(new_n934_));
  AOI211_X1 g733(.A(new_n636_), .B(new_n854_), .C1(new_n859_), .C2(new_n851_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n657_), .B1(new_n936_), .B2(new_n843_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n866_), .B(new_n938_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n756_), .B(new_n933_), .C1(new_n937_), .C2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(KEYINPUT125), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n868_), .A2(new_n942_), .A3(new_n756_), .A4(new_n933_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944_), .B2(new_n608_), .ZN(new_n945_));
  AOI211_X1 g744(.A(new_n319_), .B(new_n609_), .C1(new_n941_), .C2(new_n943_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1352gat));
  NOR2_X1   g746(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n865_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n944_), .B2(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n950_), .ZN(new_n952_));
  AOI211_X1 g751(.A(new_n952_), .B(new_n948_), .C1(new_n941_), .C2(new_n943_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1353gat));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n658_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(KEYINPUT127), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n956_), .B1(new_n944_), .B2(new_n959_), .ZN(new_n960_));
  AOI211_X1 g759(.A(new_n955_), .B(new_n958_), .C1(new_n941_), .C2(new_n943_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1354gat));
  INV_X1    g761(.A(G218gat), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n944_), .A2(new_n963_), .A3(new_n636_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n703_), .B1(new_n941_), .B2(new_n943_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n964_), .B1(new_n963_), .B2(new_n965_), .ZN(G1355gat));
endmodule


