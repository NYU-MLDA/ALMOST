//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_;
  XOR2_X1   g000(.A(G64gat), .B(G92gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT20), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT92), .B(G197gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n210_), .B2(G204gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(G197gat), .B2(G204gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(new_n210_), .B2(G204gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT93), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT93), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n219_), .B(new_n216_), .C1(new_n210_), .C2(G204gat), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n212_), .B1(new_n211_), .B2(KEYINPUT21), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n215_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G183gat), .ZN(new_n224_));
  INV_X1    g023(.A(G190gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT23), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT84), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(G183gat), .A3(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n230_), .B(KEYINPUT23), .C1(new_n224_), .C2(new_n225_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n224_), .A2(new_n225_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G169gat), .ZN(new_n235_));
  INV_X1    g034(.A(G176gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n242_));
  INV_X1    g041(.A(G169gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n236_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n244_), .A2(new_n245_), .B1(KEYINPUT24), .B2(new_n238_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(KEYINPUT24), .A3(new_n245_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT26), .B(G190gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT25), .B(G183gat), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n250_), .A2(new_n251_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n241_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n208_), .B1(new_n223_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT96), .Z(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT19), .Z(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n222_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n218_), .A2(new_n220_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n260_), .A2(new_n261_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT26), .B(G190gat), .Z(new_n263_));
  INV_X1    g062(.A(KEYINPUT81), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT82), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT81), .B1(new_n267_), .B2(G190gat), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n265_), .A2(new_n266_), .A3(new_n251_), .A4(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n251_), .B(new_n268_), .C1(new_n250_), .C2(KEYINPUT81), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT82), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n229_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(KEYINPUT84), .B2(new_n226_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n248_), .A2(new_n247_), .B1(new_n274_), .B2(new_n231_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n226_), .A2(new_n229_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n277_), .A2(new_n233_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(new_n239_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n262_), .A2(new_n276_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n255_), .A2(new_n259_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n223_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n240_), .A2(new_n234_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n208_), .B1(new_n262_), .B2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n259_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n207_), .B1(new_n283_), .B2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n284_), .A2(new_n223_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT20), .B1(new_n262_), .B2(new_n286_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n258_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n285_), .A2(new_n287_), .A3(new_n259_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n206_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(KEYINPUT27), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT99), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n285_), .A2(new_n287_), .A3(new_n259_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n259_), .B1(new_n255_), .B2(new_n281_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n207_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n294_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n295_), .A2(new_n296_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT91), .B(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT90), .B(G228gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT94), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n305_), .B1(new_n262_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G78gat), .B(G106gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OR4_X1    g108(.A1(KEYINPUT87), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT86), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n317_));
  INV_X1    g116(.A(G141gat), .ZN(new_n318_));
  INV_X1    g117(.A(G148gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(KEYINPUT87), .B2(KEYINPUT3), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n310_), .A2(new_n316_), .A3(new_n317_), .A4(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G155gat), .B(G162gat), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT1), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n312_), .A2(new_n314_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n320_), .A4(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n309_), .B1(new_n223_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n324_), .B2(new_n329_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n262_), .A2(new_n308_), .A3(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n307_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n308_), .B1(new_n262_), .B2(new_n334_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n223_), .A2(new_n309_), .A3(new_n331_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n223_), .A2(KEYINPUT94), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .A4(new_n305_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(KEYINPUT89), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT95), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT95), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n336_), .A2(new_n343_), .A3(new_n340_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G22gat), .B(G50gat), .Z(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n330_), .B2(KEYINPUT29), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT88), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n324_), .A2(new_n348_), .A3(new_n329_), .A4(new_n333_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n346_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n345_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT88), .ZN(new_n354_));
  INV_X1    g153(.A(new_n345_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n346_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n342_), .A2(new_n344_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(new_n357_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n341_), .A3(KEYINPUT95), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT98), .B(KEYINPUT0), .Z(new_n363_));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G57gat), .B(G85gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G127gat), .B(G134gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n369_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(KEYINPUT85), .A3(new_n371_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n330_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n324_), .A2(new_n372_), .A3(new_n329_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(KEYINPUT4), .ZN(new_n381_));
  INV_X1    g180(.A(new_n375_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT85), .B1(new_n370_), .B2(new_n371_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT4), .B1(new_n384_), .B2(new_n330_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n367_), .B(new_n380_), .C1(new_n387_), .C2(new_n379_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n367_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n391_), .A2(new_n385_), .A3(new_n379_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n380_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n389_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n374_), .A2(new_n375_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT31), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n397_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G43gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT30), .B1(new_n276_), .B2(new_n280_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT30), .ZN(new_n404_));
  AOI211_X1 g203(.A(new_n404_), .B(new_n279_), .C1(new_n272_), .C2(new_n275_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n248_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n232_), .B1(new_n409_), .B2(new_n246_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n271_), .B2(new_n269_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n404_), .B1(new_n411_), .B2(new_n279_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n276_), .A2(KEYINPUT30), .A3(new_n280_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n401_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n408_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n408_), .B1(new_n406_), .B2(new_n414_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n400_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n406_), .A2(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n407_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n397_), .B(new_n398_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n415_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n395_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n289_), .A2(KEYINPUT99), .A3(KEYINPUT27), .A4(new_n294_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n302_), .A2(new_n362_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT100), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n294_), .A2(KEYINPUT27), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n262_), .B1(new_n280_), .B2(new_n276_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT20), .B1(new_n223_), .B2(new_n254_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n258_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n206_), .B1(new_n431_), .B2(new_n282_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n296_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n300_), .A2(new_n301_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n424_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n435_), .A2(KEYINPUT100), .A3(new_n362_), .A4(new_n423_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n427_), .A2(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(KEYINPUT33), .B(new_n389_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n438_), .A2(new_n294_), .A3(new_n299_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n367_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n387_), .B2(new_n379_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n394_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n431_), .B2(new_n282_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n297_), .A2(new_n298_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n439_), .A2(new_n443_), .B1(new_n447_), .B2(new_n395_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n359_), .A2(new_n361_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n433_), .A2(new_n434_), .A3(new_n424_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n395_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n359_), .A2(new_n451_), .A3(new_n361_), .ZN(new_n452_));
  OAI22_X1  g251(.A1(new_n448_), .A2(new_n449_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n418_), .A2(new_n422_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n437_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G230gat), .ZN(new_n457_));
  INV_X1    g256(.A(G233gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G64gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(G57gat), .ZN(new_n461_));
  INV_X1    g260(.A(G57gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G64gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT11), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G71gat), .B(G78gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT69), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(G71gat), .A2(G78gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G71gat), .A2(G78gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT69), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G57gat), .B(G64gat), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n469_), .B(new_n470_), .C1(new_n471_), .C2(KEYINPUT11), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n466_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(KEYINPUT11), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n474_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n466_), .A2(new_n476_), .A3(new_n472_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n479_));
  INV_X1    g278(.A(G99gat), .ZN(new_n480_));
  INV_X1    g279(.A(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(KEYINPUT66), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n483_), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n479_), .B1(new_n486_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n490_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(new_n487_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n493_), .A2(new_n495_), .A3(KEYINPUT67), .A4(new_n489_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n492_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504_));
  OR2_X1    g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n497_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n497_), .A2(new_n504_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT65), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT9), .B1(new_n498_), .B2(new_n499_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT65), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n507_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n488_), .A2(new_n490_), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT10), .B(G99gat), .Z(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT64), .B(G106gat), .Z(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT68), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT68), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT6), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n525_), .A2(new_n493_), .A3(new_n489_), .A4(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n500_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(new_n502_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n513_), .A2(new_n517_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n478_), .A2(new_n503_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT70), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n478_), .A2(new_n503_), .A3(KEYINPUT70), .A4(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n478_), .B1(new_n503_), .B2(new_n530_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n459_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n459_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n466_), .A2(new_n476_), .A3(new_n472_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n476_), .B1(new_n466_), .B2(new_n472_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n493_), .A2(new_n495_), .A3(new_n489_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n528_), .B1(new_n544_), .B2(new_n479_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT8), .B1(new_n545_), .B2(new_n496_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n506_), .A2(KEYINPUT65), .A3(new_n508_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n511_), .B1(new_n510_), .B2(new_n507_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n517_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n527_), .A2(new_n529_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n543_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT12), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT12), .B1(new_n552_), .B2(new_n553_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n540_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n537_), .A2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT73), .B(KEYINPUT5), .Z(new_n558_));
  XNOR2_X1  g357(.A(G120gat), .B(G148gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G176gat), .B(G204gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT72), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n557_), .B(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT75), .B(G1gat), .ZN(new_n567_));
  INV_X1    g366(.A(G8gat), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT14), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G1gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n570_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n573_), .A2(new_n568_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(new_n571_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(G1gat), .ZN(new_n577_));
  AOI21_X1  g376(.A(G8gat), .B1(new_n577_), .B2(new_n572_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n568_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(G8gat), .A3(new_n572_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(G231gat), .A3(G233gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n478_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n581_), .A2(new_n585_), .A3(new_n543_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT76), .A3(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT16), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G183gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G211gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n589_), .B(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(KEYINPUT17), .ZN(new_n596_));
  INV_X1    g395(.A(new_n587_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n588_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G169gat), .B(G197gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT79), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  XNOR2_X1  g404(.A(G29gat), .B(G36gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G43gat), .B(G50gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT77), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n584_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n608_), .B(KEYINPUT15), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT78), .B1(new_n614_), .B2(new_n584_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT78), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n579_), .A2(new_n616_), .A3(new_n613_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n612_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n609_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n579_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n611_), .B1(new_n620_), .B2(new_n610_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n605_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n610_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n611_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n605_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n615_), .A2(new_n617_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n625_), .B(new_n626_), .C1(new_n627_), .C2(new_n612_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT80), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT80), .B(new_n605_), .C1(new_n618_), .C2(new_n621_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n566_), .A2(new_n600_), .A3(new_n601_), .A4(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n546_), .A2(new_n551_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n608_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n613_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT34), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT35), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n638_), .A2(KEYINPUT74), .A3(new_n639_), .A4(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(KEYINPUT35), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G190gat), .B(G218gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(KEYINPUT36), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n648_), .B(KEYINPUT36), .Z(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n645_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n636_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n650_), .B(KEYINPUT37), .C1(new_n645_), .C2(new_n653_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n456_), .A2(new_n635_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n395_), .A3(new_n567_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT102), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT102), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n634_), .B(KEYINPUT103), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n651_), .A2(new_n654_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n668_), .A2(new_n456_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n451_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n663_), .A2(KEYINPUT38), .A3(new_n664_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n667_), .A2(new_n673_), .A3(new_n674_), .ZN(G1324gat));
  NAND3_X1  g474(.A1(new_n661_), .A2(new_n568_), .A3(new_n450_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n668_), .A2(new_n450_), .A3(new_n456_), .A4(new_n670_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n677_), .A2(new_n678_), .A3(G8gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n677_), .B2(G8gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT104), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n676_), .B(new_n683_), .C1(new_n680_), .C2(new_n679_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n682_), .A2(KEYINPUT40), .A3(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n454_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n671_), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT41), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n690_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n659_), .B2(new_n694_), .ZN(G1326gat));
  INV_X1    g494(.A(G22gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n671_), .B2(new_n449_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT42), .Z(new_n698_));
  NOR2_X1   g497(.A1(new_n362_), .A2(G22gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT105), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n659_), .B2(new_n700_), .ZN(G1327gat));
  AOI22_X1  g500(.A1(new_n427_), .A2(new_n436_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n702_), .A2(new_n600_), .A3(new_n670_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n566_), .A2(new_n601_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n632_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n395_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n600_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n702_), .B2(new_n658_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n456_), .A2(new_n711_), .A3(new_n657_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT44), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n714_), .A2(G29gat), .A3(new_n395_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n709_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n711_), .B1(new_n456_), .B2(new_n657_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT43), .B(new_n658_), .C1(new_n437_), .C2(new_n455_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n707_), .B1(new_n715_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT106), .ZN(G1328gat));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n706_), .A2(new_n724_), .A3(new_n450_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT45), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n435_), .B1(new_n713_), .B2(KEYINPUT44), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n721_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n729_), .B2(G36gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT107), .B(new_n724_), .C1(new_n728_), .C2(new_n721_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(KEYINPUT46), .B(new_n726_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1329gat));
  NAND3_X1  g535(.A1(new_n714_), .A2(G43gat), .A3(new_n691_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n721_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n706_), .A2(new_n691_), .ZN(new_n739_));
  OAI22_X1  g538(.A1(new_n737_), .A2(new_n738_), .B1(G43gat), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g540(.A1(new_n714_), .A2(G50gat), .A3(new_n449_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n706_), .A2(new_n449_), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n742_), .A2(new_n738_), .B1(G50gat), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT108), .ZN(G1331gat));
  INV_X1    g544(.A(new_n704_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n702_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n655_), .A2(new_n632_), .A3(new_n600_), .A4(new_n656_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n462_), .B1(new_n750_), .B2(new_n451_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT109), .Z(new_n752_));
  AND4_X1   g551(.A1(new_n632_), .A2(new_n747_), .A3(new_n600_), .A4(new_n670_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n451_), .A2(new_n462_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(G1332gat));
  AOI21_X1  g554(.A(new_n460_), .B1(new_n753_), .B2(new_n450_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT48), .Z(new_n757_));
  INV_X1    g556(.A(new_n750_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n460_), .A3(new_n450_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n753_), .B2(new_n691_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT49), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n761_), .A3(new_n691_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1334gat));
  INV_X1    g564(.A(G78gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n753_), .B2(new_n449_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT50), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n758_), .A2(new_n766_), .A3(new_n449_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n746_), .A2(new_n633_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n703_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n395_), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT110), .Z(new_n775_));
  NAND2_X1  g574(.A1(new_n710_), .A2(new_n712_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n771_), .A2(new_n708_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(G85gat), .A3(new_n395_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n775_), .A2(new_n781_), .ZN(G1336gat));
  AOI21_X1  g581(.A(G92gat), .B1(new_n773_), .B2(new_n450_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n450_), .A2(G92gat), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT111), .Z(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n780_), .B2(new_n785_), .ZN(G1337gat));
  NAND2_X1  g585(.A1(new_n780_), .A2(new_n691_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n691_), .A2(new_n515_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n787_), .A2(G99gat), .B1(new_n773_), .B2(new_n788_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g589(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n776_), .A2(new_n449_), .A3(new_n778_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(G106gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(G106gat), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n773_), .A2(new_n449_), .A3(new_n516_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n791_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n791_), .B(new_n797_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  NOR4_X1   g600(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .A4(new_n454_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n537_), .A2(new_n556_), .A3(new_n563_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n630_), .A2(new_n631_), .A3(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n554_), .A2(new_n555_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n459_), .B1(new_n807_), .B2(new_n535_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT12), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n536_), .B2(KEYINPUT71), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT12), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n539_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT55), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n556_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n808_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n562_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT56), .B1(new_n816_), .B2(new_n562_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n806_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n624_), .B1(new_n620_), .B2(new_n610_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n626_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n615_), .A2(new_n617_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n610_), .A3(new_n624_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n821_), .A2(new_n820_), .A3(new_n626_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n628_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n565_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n669_), .B1(new_n819_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n804_), .B1(new_n830_), .B2(KEYINPUT116), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n630_), .A2(new_n631_), .A3(new_n805_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n535_), .B1(new_n811_), .B2(new_n810_), .ZN(new_n833_));
  OAI22_X1  g632(.A1(new_n833_), .A2(new_n538_), .B1(new_n812_), .B2(KEYINPUT55), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n556_), .A2(new_n814_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n562_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n562_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n832_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n670_), .B1(new_n840_), .B2(new_n828_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n831_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n805_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n827_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT58), .B(new_n846_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n657_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n838_), .A2(new_n839_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n846_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT118), .B1(new_n848_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n846_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n849_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n657_), .A4(new_n847_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n830_), .A2(KEYINPUT57), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n853_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n708_), .B1(new_n844_), .B2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n704_), .B2(new_n748_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT114), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n865_), .B(new_n862_), .C1(new_n704_), .C2(new_n748_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n746_), .A2(new_n749_), .A3(new_n861_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n803_), .B1(new_n860_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(G113gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n633_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n803_), .A2(KEYINPUT119), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT59), .B1(new_n803_), .B2(KEYINPUT119), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n841_), .A2(new_n842_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n830_), .A2(KEYINPUT116), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n804_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n848_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n877_), .A2(new_n855_), .B1(new_n830_), .B2(KEYINPUT57), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n600_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n868_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n872_), .B(new_n873_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n869_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT120), .B(new_n881_), .C1(new_n869_), .C2(new_n882_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n632_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n871_), .B1(new_n887_), .B2(new_n870_), .ZN(G1340gat));
  NOR2_X1   g687(.A1(new_n746_), .A2(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n869_), .B1(KEYINPUT60), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n704_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G120gat), .B1(new_n891_), .B2(new_n883_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(KEYINPUT60), .B2(new_n890_), .ZN(G1341gat));
  AOI211_X1 g692(.A(new_n708_), .B(new_n803_), .C1(new_n860_), .C2(new_n868_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT121), .B1(new_n894_), .B2(G127gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n869_), .A2(new_n600_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897_));
  INV_X1    g696(.A(G127gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n885_), .A2(new_n886_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT122), .B(G127gat), .Z(new_n902_));
  NOR2_X1   g701(.A1(new_n708_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1342gat));
  INV_X1    g703(.A(G134gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n869_), .A2(new_n905_), .A3(new_n669_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n658_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n905_), .ZN(G1343gat));
  NAND2_X1  g707(.A1(new_n860_), .A2(new_n868_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n691_), .A2(new_n451_), .A3(new_n362_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n435_), .A3(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n632_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n318_), .ZN(G1344gat));
  NOR2_X1   g712(.A1(new_n911_), .A2(new_n746_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n319_), .ZN(G1345gat));
  NOR2_X1   g714(.A1(new_n911_), .A2(new_n708_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT61), .B(G155gat), .Z(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  OAI21_X1  g717(.A(G162gat), .B1(new_n911_), .B2(new_n658_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n670_), .A2(G162gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n911_), .B2(new_n920_), .ZN(G1347gat));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n450_), .A2(new_n423_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n449_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n633_), .B(new_n924_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n922_), .B1(new_n926_), .B2(new_n243_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(KEYINPUT62), .A3(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n235_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n929_), .B(new_n930_), .C1(KEYINPUT62), .C2(new_n927_), .ZN(G1348gat));
  OR2_X1    g730(.A1(new_n879_), .A2(new_n880_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n924_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n236_), .B1(new_n933_), .B2(new_n746_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n746_), .A2(new_n236_), .A3(new_n923_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n909_), .A2(new_n362_), .A3(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n934_), .A2(KEYINPUT124), .A3(new_n936_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1349gat));
  INV_X1    g740(.A(new_n933_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n708_), .A2(new_n251_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n708_), .A2(new_n923_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n909_), .A2(new_n362_), .A3(new_n944_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n942_), .A2(new_n943_), .B1(new_n224_), .B2(new_n945_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n933_), .B2(new_n658_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n669_), .A2(new_n250_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(KEYINPUT125), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n932_), .A2(new_n924_), .A3(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n947_), .A2(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n947_), .A2(KEYINPUT126), .A3(new_n950_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1351gat));
  NOR3_X1   g754(.A1(new_n435_), .A2(new_n691_), .A3(new_n452_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n909_), .A2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n633_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g759(.A1(new_n957_), .A2(new_n746_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n962_), .ZN(G1353gat));
  NOR2_X1   g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  AND2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  NOR4_X1   g764(.A1(new_n957_), .A2(new_n708_), .A3(new_n964_), .A4(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n958_), .A2(new_n600_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n967_), .B2(new_n964_), .ZN(G1354gat));
  OR3_X1    g767(.A1(new_n957_), .A2(G218gat), .A3(new_n670_), .ZN(new_n969_));
  OAI21_X1  g768(.A(G218gat), .B1(new_n957_), .B2(new_n658_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1355gat));
endmodule


